VERSION 5.3 ;
   NAMESCASESENSITIVE ON ;
   NOWIREEXTENSIONATPIN ON ;
   DIVIDERCHAR "/" ;
   BUSBITCHARS "[]" ;
UNITS
   DATABASE MICRONS 1000 ;
END UNITS

MACRO single_generate
   CLASS BLOCK ;
   FOREIGN single_generate ;
   ORIGIN 3.5000 1.0000 ;
   SIZE 55.0000 BY 27.3000 ;
   PIN vdd
      DIRECTION INOUT ;
      PORT
         LAYER M1 ;
	    RECT 2.8000 1.6000 3.6000 9.0000 ;
	    RECT 7.6000 1.6000 8.4000 9.0000 ;
	    RECT 12.4000 1.6000 13.2000 6.2000 ;
	    RECT 20.4000 1.6000 21.2000 10.2000 ;
	    RECT 25.2000 1.6000 26.0000 10.2000 ;
	    RECT 36.4000 1.6000 37.2000 6.2000 ;
	    RECT 39.6000 1.6000 40.4000 9.8000 ;
	    RECT 44.4000 1.6000 45.2000 9.0000 ;
	    RECT 0.4000 0.4000 47.6000 1.6000 ;
         LAYER M2 ;
	    RECT 13.8000 1.4000 15.0000 1.6000 ;
	    RECT 11.5000 0.6000 17.3000 1.4000 ;
	    RECT 13.8000 0.4000 15.0000 0.6000 ;
         LAYER M3 ;
	    RECT 11.4000 0.4000 17.4000 1.6000 ;
         LAYER M4 ;
	    RECT 11.2000 -1.0000 17.6000 21.6000 ;
      END
   END vdd
   PIN gnd
      DIRECTION INOUT ;
      PORT
         LAYER M1 ;
	    RECT 0.4000 20.4000 47.6000 21.6000 ;
	    RECT 2.8000 15.8000 3.6000 20.4000 ;
	    RECT 7.6000 15.8000 8.4000 20.4000 ;
	    RECT 12.4000 17.8000 13.2000 20.4000 ;
	    RECT 20.4000 17.8000 21.2000 20.4000 ;
	    RECT 23.6000 17.8000 24.4000 20.4000 ;
	    RECT 25.2000 17.8000 26.0000 20.4000 ;
	    RECT 28.4000 17.8000 29.2000 20.4000 ;
	    RECT 39.0000 16.0000 39.8000 20.4000 ;
	    RECT 44.4000 15.8000 45.2000 20.4000 ;
         LAYER M2 ;
	    RECT 31.4000 21.4000 32.6000 21.6000 ;
	    RECT 29.1000 20.6000 34.9000 21.4000 ;
	    RECT 31.4000 20.4000 32.6000 20.6000 ;
         LAYER M3 ;
	    RECT 29.0000 20.4000 35.0000 21.6000 ;
         LAYER M4 ;
	    RECT 28.8000 -1.0000 35.2000 21.6000 ;
      END
   END gnd
   PIN g
      DIRECTION INOUT ;
      PORT
         LAYER M1 ;
	    RECT 46.0000 14.3000 46.8000 19.8000 ;
	    RECT 47.6000 14.3000 48.4000 14.4000 ;
	    RECT 46.0000 13.7000 48.4000 14.3000 ;
	    RECT 46.0000 12.4000 46.8000 13.7000 ;
	    RECT 47.6000 13.6000 48.4000 13.7000 ;
	    RECT 46.2000 10.2000 46.8000 12.4000 ;
	    RECT 46.0000 2.2000 46.8000 10.2000 ;
         LAYER M2 ;
	    RECT 47.6000 13.6000 48.4000 14.4000 ;
	    RECT 47.7000 12.4000 48.3000 13.6000 ;
	    RECT 47.6000 11.6000 48.4000 12.4000 ;
         LAYER M3 ;
	    RECT 47.6000 12.3000 48.4000 12.4000 ;
	    RECT 47.6000 11.7000 51.5000 12.3000 ;
	    RECT 47.6000 11.6000 48.4000 11.7000 ;
      END
   END g
   PIN h
      DIRECTION INOUT ;
      PORT
         LAYER M1 ;
	    RECT 1.2000 12.4000 2.0000 19.8000 ;
	    RECT 1.2000 10.2000 1.8000 12.4000 ;
	    RECT 1.2000 2.2000 2.0000 10.2000 ;
         LAYER M2 ;
	    RECT 1.2000 15.6000 2.0000 16.4000 ;
         LAYER M3 ;
	    RECT 1.2000 16.3000 2.0000 16.4000 ;
	    RECT -3.5000 15.7000 2.0000 16.3000 ;
	    RECT 1.2000 15.6000 2.0000 15.7000 ;
      END
   END h
   PIN p
      DIRECTION INOUT ;
      PORT
         LAYER M1 ;
	    RECT 6.0000 12.4000 6.8000 19.8000 ;
	    RECT 6.0000 10.2000 6.6000 12.4000 ;
	    RECT 6.0000 2.2000 6.8000 10.2000 ;
         LAYER M2 ;
	    RECT 6.0000 13.6000 6.8000 14.4000 ;
         LAYER M3 ;
	    RECT 6.0000 14.3000 6.8000 14.4000 ;
	    RECT -3.5000 13.7000 6.8000 14.3000 ;
	    RECT -3.5000 11.7000 -2.9000 13.7000 ;
	    RECT 6.0000 13.6000 6.8000 13.7000 ;
      END
   END p
   PIN x
      DIRECTION INOUT ;
      PORT
         LAYER M1 ;
	    RECT 38.4000 13.8000 39.2000 14.0000 ;
	    RECT 38.2000 13.2000 39.2000 13.8000 ;
	    RECT 38.2000 12.4000 38.8000 13.2000 ;
	    RECT 28.4000 12.3000 29.2000 12.4000 ;
	    RECT 30.0000 12.3000 30.8000 12.4000 ;
	    RECT 28.4000 11.7000 30.8000 12.3000 ;
	    RECT 28.4000 10.8000 29.2000 11.7000 ;
	    RECT 30.0000 11.6000 30.8000 11.7000 ;
	    RECT 38.0000 11.6000 38.8000 12.4000 ;
         LAYER M2 ;
	    RECT 30.0000 15.6000 30.8000 16.4000 ;
	    RECT 38.0000 15.6000 38.8000 16.4000 ;
	    RECT 30.1000 12.4000 30.7000 15.6000 ;
	    RECT 38.1000 12.4000 38.7000 15.6000 ;
	    RECT 30.0000 11.6000 30.8000 12.4000 ;
	    RECT 38.0000 11.6000 38.8000 12.4000 ;
         LAYER M3 ;
	    RECT 30.0000 16.3000 30.8000 16.4000 ;
	    RECT 38.0000 16.3000 38.8000 16.4000 ;
	    RECT 30.0000 15.7000 51.5000 16.3000 ;
	    RECT 30.0000 15.6000 30.8000 15.7000 ;
	    RECT 38.0000 15.6000 38.8000 15.7000 ;
      END
   END x
   PIN y
      DIRECTION INOUT ;
      PORT
         LAYER M1 ;
	    RECT 25.2000 15.6000 26.0000 17.2000 ;
	    RECT 28.4000 14.3000 29.2000 14.4000 ;
	    RECT 36.4000 14.3000 37.2000 14.4000 ;
	    RECT 28.4000 13.7000 37.2000 14.3000 ;
	    RECT 28.4000 13.6000 29.2000 13.7000 ;
	    RECT 36.4000 12.8000 37.2000 13.7000 ;
         LAYER M2 ;
	    RECT 25.3000 18.4000 25.9000 26.3000 ;
	    RECT 25.2000 17.6000 26.0000 18.4000 ;
	    RECT 28.4000 17.6000 29.2000 18.4000 ;
	    RECT 25.3000 16.4000 25.9000 17.6000 ;
	    RECT 25.2000 15.6000 26.0000 16.4000 ;
	    RECT 28.5000 14.4000 29.1000 17.6000 ;
	    RECT 28.4000 13.6000 29.2000 14.4000 ;
         LAYER M3 ;
	    RECT 25.2000 18.3000 26.0000 18.4000 ;
	    RECT 28.4000 18.3000 29.2000 18.4000 ;
	    RECT 25.2000 17.7000 29.2000 18.3000 ;
	    RECT 25.2000 17.6000 26.0000 17.7000 ;
	    RECT 28.4000 17.6000 29.2000 17.7000 ;
      END
   END y
   OBS
         LAYER M1 ;
	    RECT 4.4000 15.2000 5.2000 19.8000 ;
	    RECT 9.2000 15.2000 10.0000 19.8000 ;
	    RECT 3.0000 14.6000 5.2000 15.2000 ;
	    RECT 7.8000 14.6000 10.0000 15.2000 ;
	    RECT 3.0000 11.6000 3.6000 14.6000 ;
	    RECT 4.4000 11.6000 5.2000 13.2000 ;
	    RECT 7.8000 11.6000 8.4000 14.6000 ;
	    RECT 9.2000 12.3000 10.0000 13.2000 ;
	    RECT 10.8000 12.3000 11.6000 19.8000 ;
	    RECT 22.0000 17.8000 22.8000 19.8000 ;
	    RECT 26.8000 17.8000 27.6000 19.8000 ;
	    RECT 12.4000 16.3000 13.2000 17.2000 ;
	    RECT 20.4000 16.3000 21.2000 17.2000 ;
	    RECT 12.4000 15.7000 21.2000 16.3000 ;
	    RECT 12.4000 15.6000 13.2000 15.7000 ;
	    RECT 20.4000 15.6000 21.2000 15.7000 ;
	    RECT 22.2000 14.4000 22.8000 17.8000 ;
	    RECT 27.0000 16.4000 27.6000 17.8000 ;
	    RECT 26.8000 15.6000 27.6000 16.4000 ;
	    RECT 36.4000 15.8000 37.2000 19.8000 ;
	    RECT 40.6000 16.8000 41.4000 19.8000 ;
	    RECT 40.6000 15.8000 42.0000 16.8000 ;
	    RECT 27.0000 14.4000 27.6000 15.6000 ;
	    RECT 36.6000 15.6000 37.2000 15.8000 ;
	    RECT 36.6000 15.2000 38.4000 15.6000 ;
	    RECT 36.6000 15.0000 40.8000 15.2000 ;
	    RECT 37.8000 14.6000 40.8000 15.0000 ;
	    RECT 22.0000 13.6000 22.8000 14.4000 ;
	    RECT 26.8000 13.6000 27.6000 14.4000 ;
	    RECT 9.2000 11.7000 11.6000 12.3000 ;
	    RECT 9.2000 11.6000 10.0000 11.7000 ;
	    RECT 2.4000 10.8000 3.6000 11.6000 ;
	    RECT 7.2000 10.8000 8.4000 11.6000 ;
	    RECT 3.0000 10.2000 3.6000 10.8000 ;
	    RECT 7.8000 10.2000 8.4000 10.8000 ;
	    RECT 3.0000 9.6000 5.2000 10.2000 ;
	    RECT 7.8000 9.6000 10.0000 10.2000 ;
	    RECT 4.4000 2.2000 5.2000 9.6000 ;
	    RECT 9.2000 2.2000 10.0000 9.6000 ;
	    RECT 10.8000 2.2000 11.6000 11.7000 ;
	    RECT 12.4000 12.3000 13.2000 12.4000 ;
	    RECT 22.2000 12.3000 22.8000 13.6000 ;
	    RECT 12.4000 11.7000 22.8000 12.3000 ;
	    RECT 12.4000 11.6000 13.2000 11.7000 ;
	    RECT 22.2000 10.2000 22.8000 11.7000 ;
	    RECT 23.6000 10.8000 24.4000 12.4000 ;
	    RECT 27.0000 10.2000 27.6000 13.6000 ;
	    RECT 40.0000 14.4000 40.8000 14.6000 ;
	    RECT 40.0000 11.0000 40.6000 14.4000 ;
	    RECT 41.4000 12.4000 42.0000 15.8000 ;
	    RECT 42.8000 15.2000 43.6000 19.8000 ;
	    RECT 42.8000 14.6000 45.0000 15.2000 ;
	    RECT 41.2000 12.3000 42.0000 12.4000 ;
	    RECT 42.8000 12.3000 43.6000 13.2000 ;
	    RECT 41.2000 11.7000 43.6000 12.3000 ;
	    RECT 41.2000 11.6000 42.0000 11.7000 ;
	    RECT 42.8000 11.6000 43.6000 11.7000 ;
	    RECT 44.4000 11.6000 45.0000 14.6000 ;
	    RECT 38.2000 10.4000 40.6000 11.0000 ;
	    RECT 22.0000 9.4000 23.8000 10.2000 ;
	    RECT 26.8000 9.4000 28.6000 10.2000 ;
	    RECT 23.0000 2.2000 23.8000 9.4000 ;
	    RECT 27.8000 2.2000 28.6000 9.4000 ;
	    RECT 38.2000 6.2000 38.8000 10.4000 ;
	    RECT 41.4000 10.2000 42.0000 11.6000 ;
	    RECT 44.4000 10.8000 45.6000 11.6000 ;
	    RECT 44.4000 10.2000 45.0000 10.8000 ;
	    RECT 38.0000 2.2000 38.8000 6.2000 ;
	    RECT 41.2000 2.2000 42.0000 10.2000 ;
	    RECT 42.8000 9.6000 45.0000 10.2000 ;
	    RECT 42.8000 2.2000 43.6000 9.6000 ;
         LAYER M2 ;
	    RECT 20.4000 15.6000 21.2000 16.4000 ;
	    RECT 26.8000 15.6000 27.6000 16.4000 ;
	    RECT 4.4000 11.6000 5.2000 12.4000 ;
	    RECT 12.4000 11.6000 13.2000 12.4000 ;
	    RECT 23.6000 11.6000 24.4000 12.4000 ;
	    RECT 41.2000 11.6000 42.0000 12.4000 ;
         LAYER M3 ;
	    RECT 20.4000 16.3000 21.2000 16.4000 ;
	    RECT 26.8000 16.3000 27.6000 16.4000 ;
	    RECT 20.4000 15.7000 27.6000 16.3000 ;
	    RECT 20.4000 15.6000 21.2000 15.7000 ;
	    RECT 26.8000 15.6000 27.6000 15.7000 ;
	    RECT 4.4000 12.3000 5.2000 12.4000 ;
	    RECT 12.4000 12.3000 13.2000 12.4000 ;
	    RECT 4.4000 11.7000 13.2000 12.3000 ;
	    RECT 4.4000 11.6000 5.2000 11.7000 ;
	    RECT 12.4000 11.6000 13.2000 11.7000 ;
	    RECT 23.6000 12.3000 24.4000 12.4000 ;
	    RECT 41.2000 12.3000 42.0000 12.4000 ;
	    RECT 23.6000 11.7000 42.0000 12.3000 ;
	    RECT 23.6000 11.6000 24.4000 11.7000 ;
	    RECT 41.2000 11.6000 42.0000 11.7000 ;
   END
END single_generate
