magic
tech scmos
timestamp 1592523792
<< metal1 >>
rect 181 107 187 108
rect 176 103 177 107
rect 181 103 182 107
rect 186 103 187 107
rect 191 103 192 107
rect 181 102 187 103
rect 106 78 113 81
rect 158 78 169 81
rect 102 71 105 78
rect 78 68 105 71
rect 158 68 169 71
rect 166 62 169 68
rect 22 58 30 61
rect 114 58 121 61
rect 142 58 150 61
rect 222 58 241 61
rect 254 38 262 41
rect 77 7 83 8
rect 72 3 73 7
rect 77 3 78 7
rect 82 3 83 7
rect 87 3 88 7
rect 77 2 83 3
<< m2contact >>
rect 172 103 176 107
rect 177 103 181 107
rect 182 103 186 107
rect 187 103 191 107
rect 192 103 196 107
rect 126 88 130 92
rect 102 78 106 82
rect 150 78 154 82
rect 174 78 178 82
rect 30 68 34 72
rect 214 68 218 72
rect 30 58 34 62
rect 54 58 58 62
rect 110 58 114 62
rect 150 58 154 62
rect 166 58 170 62
rect 182 58 186 62
rect 230 48 234 52
rect 6 38 10 42
rect 262 38 266 42
rect 68 3 72 7
rect 73 3 77 7
rect 78 3 82 7
rect 83 3 87 7
rect 88 3 92 7
<< metal2 >>
rect 102 138 106 142
rect 134 141 138 142
rect 126 138 138 141
rect 150 138 154 142
rect 102 82 105 138
rect 126 92 129 138
rect 150 82 153 138
rect 181 107 187 108
rect 176 103 177 107
rect 181 103 182 107
rect 186 103 187 107
rect 191 103 192 107
rect 181 102 187 103
rect 170 78 174 81
rect 30 72 33 78
rect 210 68 214 71
rect 150 62 153 68
rect 166 62 169 68
rect 26 58 30 61
rect 114 58 118 61
rect 178 58 182 61
rect 54 52 57 58
rect 230 52 233 58
rect 6 42 9 48
rect 262 42 265 48
rect 77 7 83 8
rect 72 3 73 7
rect 77 3 78 7
rect 82 3 83 7
rect 87 3 88 7
rect 77 2 83 3
<< m3contact >>
rect 172 103 176 107
rect 177 103 181 107
rect 182 103 186 107
rect 187 103 191 107
rect 192 103 196 107
rect 30 78 34 82
rect 150 78 154 82
rect 166 78 170 82
rect 150 68 154 72
rect 166 68 170 72
rect 206 68 210 72
rect 22 58 26 62
rect 118 58 122 62
rect 174 58 178 62
rect 230 58 234 62
rect 6 48 10 52
rect 54 48 58 52
rect 262 48 266 52
rect 68 3 72 7
rect 73 3 77 7
rect 78 3 82 7
rect 83 3 87 7
rect 88 3 92 7
<< metal3 >>
rect 181 107 187 108
rect 181 102 187 103
rect 34 78 150 81
rect 158 78 166 81
rect 158 71 161 78
rect 154 68 161 71
rect 170 68 206 71
rect 26 58 57 61
rect 122 58 174 61
rect 178 58 230 61
rect 54 52 57 58
rect -26 51 -22 52
rect -26 48 6 51
rect 286 51 290 52
rect 266 48 290 51
rect 77 7 83 8
rect 77 2 83 3
<< m4contact >>
rect 173 103 176 107
rect 176 103 177 107
rect 179 103 181 107
rect 181 103 182 107
rect 182 103 183 107
rect 185 103 186 107
rect 186 103 187 107
rect 187 103 189 107
rect 191 103 192 107
rect 192 103 195 107
rect 69 3 72 7
rect 72 3 73 7
rect 75 3 77 7
rect 77 3 78 7
rect 78 3 79 7
rect 81 3 82 7
rect 82 3 83 7
rect 83 3 85 7
rect 87 3 88 7
rect 88 3 91 7
<< metal4 >>
rect 181 107 187 108
rect 181 102 187 103
rect 77 7 83 8
rect 77 2 83 3
<< m5contact >>
rect 172 103 173 107
rect 173 103 176 107
rect 177 103 179 107
rect 179 103 181 107
rect 182 103 183 107
rect 183 103 185 107
rect 185 103 186 107
rect 187 103 189 107
rect 189 103 191 107
rect 192 103 195 107
rect 195 103 196 107
rect 68 3 69 7
rect 69 3 72 7
rect 73 3 75 7
rect 75 3 77 7
rect 78 3 79 7
rect 79 3 81 7
rect 81 3 82 7
rect 83 3 85 7
rect 85 3 87 7
rect 88 3 91 7
rect 91 3 92 7
<< metal5 >>
rect 181 107 187 108
rect 176 103 177 107
rect 191 103 192 107
rect 183 102 185 103
rect 77 7 83 8
rect 72 3 73 7
rect 87 3 88 7
rect 79 2 81 3
<< m6contact >>
rect 178 103 181 107
rect 181 103 182 107
rect 182 103 183 107
rect 185 103 186 107
rect 186 103 187 107
rect 187 103 190 107
rect 178 102 183 103
rect 185 102 190 103
rect 74 3 77 7
rect 77 3 78 7
rect 78 3 79 7
rect 81 3 82 7
rect 82 3 83 7
rect 83 3 86 7
rect 74 2 79 3
rect 81 2 86 3
<< metal6 >>
rect 68 7 92 107
rect 68 2 74 7
rect 79 2 81 7
rect 86 2 92 7
rect 68 -6 92 2
rect 172 102 178 107
rect 183 102 185 107
rect 190 102 196 107
rect 172 -6 196 102
use BUFX2  _11_
timestamp 1592523792
transform -1 0 28 0 -1 105
box -2 -3 26 103
use XOR2X1  _9_
timestamp 1592523792
transform 1 0 28 0 -1 105
box -2 -3 58 103
use INVX1  _6_
timestamp 1592523792
transform 1 0 108 0 -1 105
box -2 -3 18 103
use BUFX2  _10_
timestamp 1592523792
transform -1 0 148 0 -1 105
box -2 -3 26 103
use FILL  SFILL840x50
timestamp 1592523792
transform -1 0 92 0 -1 105
box -2 -3 10 103
use FILL  SFILL920x50
timestamp 1592523792
transform -1 0 100 0 -1 105
box -2 -3 10 103
use FILL  SFILL1000x50
timestamp 1592523792
transform -1 0 108 0 -1 105
box -2 -3 10 103
use INVX1  _5_
timestamp 1592523792
transform 1 0 148 0 -1 105
box -2 -3 18 103
use NOR2X1  _7_
timestamp 1592523792
transform 1 0 164 0 -1 105
box -2 -3 26 103
use NAND2X1  _8_
timestamp 1592523792
transform 1 0 212 0 -1 105
box -2 -3 26 103
use BUFX2  _12_
timestamp 1592523792
transform 1 0 236 0 -1 105
box -2 -3 26 103
use FILL  SFILL1880x50
timestamp 1592523792
transform -1 0 196 0 -1 105
box -2 -3 10 103
use FILL  SFILL1960x50
timestamp 1592523792
transform -1 0 204 0 -1 105
box -2 -3 10 103
use FILL  SFILL2040x50
timestamp 1592523792
transform -1 0 212 0 -1 105
box -2 -3 10 103
<< labels >>
flabel metal6 s 172 -6 196 0 7 FreeSans 24 270 0 0 gnd
port 0 nsew
flabel metal6 s 68 -6 92 0 7 FreeSans 24 270 0 0 vdd
port 1 nsew
flabel metal2 s 134 138 138 142 3 FreeSans 24 90 0 0 g
port 2 nsew
flabel metal3 s -26 48 -22 52 7 FreeSans 24 270 0 0 h
port 3 nsew
flabel metal3 s 286 48 290 52 3 FreeSans 24 270 0 0 p
port 4 nsew
flabel metal2 s 102 138 106 142 3 FreeSans 24 90 0 0 x
port 5 nsew
flabel metal2 s 150 138 154 142 3 FreeSans 24 90 0 0 y
port 6 nsew
<< end >>
