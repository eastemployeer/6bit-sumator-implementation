VERSION 5.3 ;
   NAMESCASESENSITIVE ON ;
   NOWIREEXTENSIONATPIN ON ;
   DIVIDERCHAR "/" ;
   BUSBITCHARS "[]" ;
UNITS
   DATABASE MICRONS 1000 ;
END UNITS

MACRO adder
   CLASS BLOCK ;
   FOREIGN adder ;
   ORIGIN 2.5500 2.1500 ;
   SIZE 69.9000 BY 36.3000 ;
   PIN gnd
      PORT
         LAYER metal1 ;
	    RECT 0.2000 30.2000 64.6000 30.8000 ;
	    RECT 1.4000 27.9000 1.8000 30.2000 ;
	    RECT 3.9000 29.9000 4.3000 30.2000 ;
	    RECT 3.8000 28.2000 4.3000 29.9000 ;
	    RECT 6.9000 28.2000 7.4000 30.2000 ;
	    RECT 9.5000 29.9000 9.9000 30.2000 ;
	    RECT 9.4000 28.2000 9.9000 29.9000 ;
	    RECT 12.5000 28.2000 13.0000 30.2000 ;
	    RECT 14.2000 28.9000 14.6000 30.2000 ;
	    RECT 15.8000 28.9000 16.2000 30.2000 ;
	    RECT 20.6000 27.9000 21.0000 30.2000 ;
	    RECT 23.1000 29.9000 23.5000 30.2000 ;
	    RECT 23.0000 28.2000 23.5000 29.9000 ;
	    RECT 26.1000 28.2000 26.6000 30.2000 ;
	    RECT 27.8000 28.9000 28.2000 30.2000 ;
	    RECT 29.4000 28.9000 29.8000 30.2000 ;
	    RECT 31.0000 28.9000 31.4000 30.2000 ;
	    RECT 31.8000 28.9000 32.2000 30.2000 ;
	    RECT 35.0000 27.9000 35.4000 30.2000 ;
	    RECT 35.8000 28.9000 36.2000 30.2000 ;
	    RECT 37.4000 28.9000 37.8000 30.2000 ;
	    RECT 39.8000 27.9000 40.2000 30.2000 ;
	    RECT 41.4000 28.9000 41.8000 30.2000 ;
	    RECT 43.0000 28.9000 43.4000 30.2000 ;
	    RECT 44.6000 28.2000 45.1000 30.2000 ;
	    RECT 47.7000 29.9000 48.1000 30.2000 ;
	    RECT 47.7000 28.2000 48.2000 29.9000 ;
	    RECT 52.6000 28.2000 53.1000 30.2000 ;
	    RECT 55.7000 29.9000 56.1000 30.2000 ;
	    RECT 55.7000 28.2000 56.2000 29.9000 ;
	    RECT 58.2000 28.9000 58.6000 30.2000 ;
	    RECT 59.8000 27.9000 60.2000 30.2000 ;
	    RECT 62.2000 27.9000 62.6000 30.2000 ;
	    RECT 1.4000 10.8000 1.9000 12.8000 ;
	    RECT 4.5000 11.1000 5.0000 12.8000 ;
	    RECT 4.5000 10.8000 4.9000 11.1000 ;
	    RECT 6.2000 10.8000 6.6000 12.1000 ;
	    RECT 7.8000 10.8000 8.2000 12.1000 ;
	    RECT 9.4000 10.8000 9.8000 12.1000 ;
	    RECT 11.0000 10.8000 11.4000 12.1000 ;
	    RECT 11.8000 10.8000 12.2000 13.1000 ;
	    RECT 15.8000 10.8000 16.2000 13.1000 ;
	    RECT 19.0000 10.8000 19.4000 12.1000 ;
	    RECT 20.6000 10.8000 21.0000 12.1000 ;
	    RECT 21.4000 10.8000 21.8000 13.1000 ;
	    RECT 23.8000 10.8000 24.2000 12.1000 ;
	    RECT 25.4000 10.8000 25.8000 13.1000 ;
	    RECT 28.6000 10.8000 29.1000 12.8000 ;
	    RECT 31.7000 11.1000 32.2000 12.8000 ;
	    RECT 31.7000 10.8000 32.1000 11.1000 ;
	    RECT 35.0000 10.8000 35.4000 13.1000 ;
	    RECT 35.8000 10.8000 36.2000 12.1000 ;
	    RECT 37.4000 10.8000 37.8000 13.1000 ;
	    RECT 41.1000 10.8000 41.5000 13.0000 ;
	    RECT 44.6000 10.8000 45.0000 13.1000 ;
	    RECT 47.0000 10.8000 47.4000 13.1000 ;
	    RECT 50.2000 10.8000 50.6000 12.1000 ;
	    RECT 51.8000 10.8000 52.2000 13.1000 ;
	    RECT 55.8000 10.8000 56.2000 13.1000 ;
	    RECT 57.4000 10.8000 57.9000 12.8000 ;
	    RECT 60.5000 11.1000 61.0000 12.8000 ;
	    RECT 60.5000 10.8000 60.9000 11.1000 ;
	    RECT 63.0000 10.8000 63.4000 13.1000 ;
	    RECT 0.2000 10.2000 64.6000 10.8000 ;
	    RECT 1.4000 7.9000 1.8000 10.2000 ;
	    RECT 3.8000 8.2000 4.3000 10.2000 ;
	    RECT 6.9000 9.9000 7.3000 10.2000 ;
	    RECT 6.9000 8.2000 7.4000 9.9000 ;
	    RECT 8.6000 7.9000 9.0000 10.2000 ;
	    RECT 12.6000 7.9000 13.0000 10.2000 ;
	    RECT 14.2000 8.9000 14.6000 10.2000 ;
	    RECT 16.3000 8.0000 16.7000 10.2000 ;
	    RECT 22.2000 7.9000 22.6000 10.2000 ;
	    RECT 24.6000 7.9000 25.0000 10.2000 ;
	    RECT 26.2000 8.9000 26.6000 10.2000 ;
	    RECT 27.8000 7.9000 28.2000 10.2000 ;
	    RECT 29.4000 8.9000 29.8000 10.2000 ;
	    RECT 31.0000 7.9000 31.4000 10.2000 ;
	    RECT 33.4000 8.9000 33.8000 10.2000 ;
	    RECT 35.0000 7.9000 35.4000 10.2000 ;
	    RECT 38.2000 8.9000 38.6000 10.2000 ;
	    RECT 39.0000 8.9000 39.4000 10.2000 ;
	    RECT 40.6000 8.9000 41.0000 10.2000 ;
	    RECT 41.4000 7.9000 41.8000 10.2000 ;
	    RECT 44.6000 8.9000 45.0000 10.2000 ;
	    RECT 48.6000 8.2000 49.1000 10.2000 ;
	    RECT 51.7000 9.9000 52.1000 10.2000 ;
	    RECT 51.7000 8.2000 52.2000 9.9000 ;
	    RECT 54.2000 8.9000 54.6000 10.2000 ;
	    RECT 55.0000 8.9000 55.4000 10.2000 ;
	    RECT 56.6000 8.9000 57.0000 10.2000 ;
	    RECT 58.3000 9.9000 58.7000 10.2000 ;
	    RECT 58.2000 8.2000 58.7000 9.9000 ;
	    RECT 61.3000 8.2000 61.8000 10.2000 ;
         LAYER metal2 ;
	    RECT 46.9000 30.7000 47.5000 30.8000 ;
	    RECT 46.0000 30.3000 48.4000 30.7000 ;
	    RECT 46.9000 30.2000 47.5000 30.3000 ;
	    RECT 46.9000 10.7000 47.5000 10.8000 ;
	    RECT 46.0000 10.3000 48.4000 10.7000 ;
	    RECT 46.9000 10.2000 47.5000 10.3000 ;
         LAYER metal3 ;
	    RECT 46.9000 30.7000 47.5000 30.8000 ;
	    RECT 46.0000 30.3000 48.4000 30.7000 ;
	    RECT 46.9000 30.2000 47.5000 30.3000 ;
	    RECT 46.9000 10.7000 47.5000 10.8000 ;
	    RECT 46.0000 10.3000 48.4000 10.7000 ;
	    RECT 46.9000 10.2000 47.5000 10.3000 ;
         LAYER metal4 ;
	    RECT 46.9000 30.7000 47.5000 30.8000 ;
	    RECT 46.0000 30.3000 48.4000 30.7000 ;
	    RECT 46.9000 30.2000 47.5000 30.3000 ;
	    RECT 46.9000 10.7000 47.5000 10.8000 ;
	    RECT 46.0000 10.3000 48.4000 10.7000 ;
	    RECT 46.9000 10.2000 47.5000 10.3000 ;
         LAYER metal5 ;
	    RECT 46.9000 30.7500 47.5000 30.8000 ;
	    RECT 46.6000 30.7000 47.8000 30.7500 ;
	    RECT 46.0000 30.3000 48.4000 30.7000 ;
	    RECT 46.6000 30.2500 47.8000 30.3000 ;
	    RECT 46.9000 30.2000 47.5000 30.2500 ;
	    RECT 46.9000 10.7500 47.5000 10.8000 ;
	    RECT 46.6000 10.7000 47.8000 10.7500 ;
	    RECT 46.0000 10.3000 48.4000 10.7000 ;
	    RECT 46.6000 10.2500 47.8000 10.3000 ;
	    RECT 46.9000 10.2000 47.5000 10.2500 ;
         LAYER metal6 ;
	    RECT 46.0000 -0.5000 48.4000 30.7500 ;
      END
   END gnd
   PIN vdd
      PORT
         LAYER metal1 ;
	    RECT 1.4000 20.8000 1.8000 24.5000 ;
	    RECT 3.8000 21.1000 4.3000 24.4000 ;
	    RECT 3.9000 20.8000 4.3000 21.1000 ;
	    RECT 6.9000 20.8000 7.4000 24.4000 ;
	    RECT 9.4000 21.1000 9.9000 24.4000 ;
	    RECT 9.5000 20.8000 9.9000 21.1000 ;
	    RECT 12.5000 20.8000 13.0000 24.4000 ;
	    RECT 14.2000 20.8000 14.6000 23.1000 ;
	    RECT 15.8000 20.8000 16.2000 23.1000 ;
	    RECT 20.6000 20.8000 21.0000 24.5000 ;
	    RECT 23.0000 21.1000 23.5000 24.4000 ;
	    RECT 23.1000 20.8000 23.5000 21.1000 ;
	    RECT 26.1000 20.8000 26.6000 24.4000 ;
	    RECT 27.8000 20.8000 28.2000 23.1000 ;
	    RECT 29.4000 20.8000 29.8000 25.1000 ;
	    RECT 31.8000 20.8000 32.2000 23.1000 ;
	    RECT 33.4000 20.8000 33.8000 23.1000 ;
	    RECT 35.0000 20.8000 35.4000 23.1000 ;
	    RECT 37.4000 20.8000 37.8000 25.1000 ;
	    RECT 38.2000 20.8000 38.6000 23.1000 ;
	    RECT 39.8000 20.8000 40.2000 23.1000 ;
	    RECT 41.4000 20.8000 41.8000 23.1000 ;
	    RECT 43.0000 20.8000 43.4000 23.1000 ;
	    RECT 44.6000 20.8000 45.1000 24.4000 ;
	    RECT 47.7000 21.1000 48.2000 24.4000 ;
	    RECT 47.7000 20.8000 48.1000 21.1000 ;
	    RECT 52.6000 20.8000 53.1000 24.4000 ;
	    RECT 55.7000 21.1000 56.2000 24.4000 ;
	    RECT 55.7000 20.8000 56.1000 21.1000 ;
	    RECT 58.2000 20.8000 58.6000 23.1000 ;
	    RECT 59.8000 20.8000 60.2000 24.5000 ;
	    RECT 62.2000 20.8000 62.6000 24.5000 ;
	    RECT 0.2000 20.2000 64.6000 20.8000 ;
	    RECT 1.4000 16.6000 1.9000 20.2000 ;
	    RECT 4.5000 19.9000 4.9000 20.2000 ;
	    RECT 4.5000 16.6000 5.0000 19.9000 ;
	    RECT 6.2000 17.9000 6.6000 20.2000 ;
	    RECT 7.8000 17.9000 8.2000 20.2000 ;
	    RECT 11.0000 15.9000 11.4000 20.2000 ;
	    RECT 11.8000 17.9000 12.2000 20.2000 ;
	    RECT 13.4000 17.9000 13.8000 20.2000 ;
	    RECT 14.2000 17.9000 14.6000 20.2000 ;
	    RECT 15.8000 17.9000 16.2000 20.2000 ;
	    RECT 20.6000 15.9000 21.0000 20.2000 ;
	    RECT 21.4000 17.9000 21.8000 20.2000 ;
	    RECT 23.0000 17.9000 23.4000 20.2000 ;
	    RECT 23.8000 17.9000 24.2000 20.2000 ;
	    RECT 25.4000 17.9000 25.8000 20.2000 ;
	    RECT 27.0000 17.9000 27.4000 20.2000 ;
	    RECT 28.6000 16.6000 29.1000 20.2000 ;
	    RECT 31.7000 19.9000 32.1000 20.2000 ;
	    RECT 31.7000 16.6000 32.2000 19.9000 ;
	    RECT 33.4000 17.9000 33.8000 20.2000 ;
	    RECT 35.0000 17.9000 35.4000 20.2000 ;
	    RECT 35.8000 17.9000 36.2000 20.2000 ;
	    RECT 37.4000 17.9000 37.8000 20.2000 ;
	    RECT 39.0000 17.9000 39.4000 20.2000 ;
	    RECT 39.8000 17.9000 40.2000 20.2000 ;
	    RECT 41.4000 16.1000 41.8000 20.2000 ;
	    RECT 43.0000 17.9000 43.4000 20.2000 ;
	    RECT 44.6000 17.9000 45.0000 20.2000 ;
	    RECT 45.4000 17.9000 45.8000 20.2000 ;
	    RECT 47.0000 17.9000 47.4000 20.2000 ;
	    RECT 50.2000 17.9000 50.6000 20.2000 ;
	    RECT 51.8000 17.9000 52.2000 20.2000 ;
	    RECT 53.4000 17.9000 53.8000 20.2000 ;
	    RECT 54.2000 17.9000 54.6000 20.2000 ;
	    RECT 55.8000 17.9000 56.2000 20.2000 ;
	    RECT 57.4000 16.6000 57.9000 20.2000 ;
	    RECT 60.5000 19.9000 60.9000 20.2000 ;
	    RECT 60.5000 16.6000 61.0000 19.9000 ;
	    RECT 63.0000 16.5000 63.4000 20.2000 ;
	    RECT 1.4000 0.8000 1.8000 4.5000 ;
	    RECT 3.8000 0.8000 4.3000 4.4000 ;
	    RECT 6.9000 1.1000 7.4000 4.4000 ;
	    RECT 6.9000 0.8000 7.3000 1.1000 ;
	    RECT 8.6000 0.8000 9.0000 3.1000 ;
	    RECT 10.2000 0.8000 10.6000 3.1000 ;
	    RECT 11.0000 0.8000 11.4000 3.1000 ;
	    RECT 12.6000 0.8000 13.0000 3.1000 ;
	    RECT 14.2000 0.8000 14.6000 3.1000 ;
	    RECT 15.0000 0.8000 15.4000 3.1000 ;
	    RECT 16.6000 0.8000 17.0000 4.9000 ;
	    RECT 20.6000 0.8000 21.0000 3.1000 ;
	    RECT 22.2000 0.8000 22.6000 3.1000 ;
	    RECT 23.0000 0.8000 23.4000 3.1000 ;
	    RECT 24.6000 0.8000 25.0000 3.1000 ;
	    RECT 26.2000 0.8000 26.6000 3.1000 ;
	    RECT 27.8000 0.8000 28.2000 4.5000 ;
	    RECT 29.4000 0.8000 29.8000 3.1000 ;
	    RECT 31.0000 0.8000 31.4000 3.1000 ;
	    RECT 32.6000 0.8000 33.0000 3.1000 ;
	    RECT 33.4000 0.8000 33.8000 3.1000 ;
	    RECT 35.0000 0.8000 35.4000 3.1000 ;
	    RECT 36.6000 0.8000 37.0000 3.1000 ;
	    RECT 38.2000 0.8000 38.6000 3.1000 ;
	    RECT 39.0000 0.8000 39.4000 5.1000 ;
	    RECT 41.4000 0.8000 41.8000 3.1000 ;
	    RECT 43.0000 0.8000 43.4000 3.1000 ;
	    RECT 44.6000 0.8000 45.0000 3.1000 ;
	    RECT 48.6000 0.8000 49.1000 4.4000 ;
	    RECT 51.7000 1.1000 52.2000 4.4000 ;
	    RECT 51.7000 0.8000 52.1000 1.1000 ;
	    RECT 54.2000 0.8000 54.6000 3.1000 ;
	    RECT 55.0000 0.8000 55.4000 5.1000 ;
	    RECT 58.2000 1.1000 58.7000 4.4000 ;
	    RECT 58.3000 0.8000 58.7000 1.1000 ;
	    RECT 61.3000 0.8000 61.8000 4.4000 ;
	    RECT 0.2000 0.2000 64.6000 0.8000 ;
         LAYER metal2 ;
	    RECT 17.3000 20.7000 17.9000 20.8000 ;
	    RECT 16.4000 20.3000 18.8000 20.7000 ;
	    RECT 17.3000 20.2000 17.9000 20.3000 ;
	    RECT 17.3000 0.7000 17.9000 0.8000 ;
	    RECT 16.4000 0.3000 18.8000 0.7000 ;
	    RECT 17.3000 0.2000 17.9000 0.3000 ;
         LAYER metal3 ;
	    RECT 17.3000 20.7000 17.9000 20.8000 ;
	    RECT 16.4000 20.3000 18.8000 20.7000 ;
	    RECT 17.3000 20.2000 17.9000 20.3000 ;
	    RECT 17.3000 0.7000 17.9000 0.8000 ;
	    RECT 16.4000 0.3000 18.8000 0.7000 ;
	    RECT 17.3000 0.2000 17.9000 0.3000 ;
         LAYER metal4 ;
	    RECT 17.3000 20.7000 17.9000 20.8000 ;
	    RECT 16.4000 20.3000 18.8000 20.7000 ;
	    RECT 17.3000 20.2000 17.9000 20.3000 ;
	    RECT 17.3000 0.7000 17.9000 0.8000 ;
	    RECT 16.4000 0.3000 18.8000 0.7000 ;
	    RECT 17.3000 0.2000 17.9000 0.3000 ;
         LAYER metal5 ;
	    RECT 17.3000 20.7500 17.9000 20.8000 ;
	    RECT 17.0000 20.7000 18.2000 20.7500 ;
	    RECT 16.4000 20.3000 18.8000 20.7000 ;
	    RECT 17.0000 20.2500 18.2000 20.3000 ;
	    RECT 17.3000 20.2000 17.9000 20.2500 ;
	    RECT 17.3000 0.7500 17.9000 0.8000 ;
	    RECT 17.0000 0.7000 18.2000 0.7500 ;
	    RECT 16.4000 0.3000 18.8000 0.7000 ;
	    RECT 17.0000 0.2500 18.2000 0.3000 ;
	    RECT 17.3000 0.2000 17.9000 0.2500 ;
         LAYER metal6 ;
	    RECT 16.4000 -0.5000 18.8000 30.7500 ;
      END
   END vdd
   PIN s[6]
      PORT
         LAYER metal1 ;
	    RECT 19.8000 26.2000 20.2000 29.9000 ;
	    RECT 19.8000 25.1000 20.1000 26.2000 ;
	    RECT 19.8000 21.1000 20.2000 25.1000 ;
         LAYER metal2 ;
	    RECT 21.4500 30.2000 21.7500 34.1500 ;
	    RECT 19.8000 29.8000 20.2000 30.2000 ;
	    RECT 21.4000 29.8000 21.8000 30.2000 ;
	    RECT 19.8500 29.2000 20.1500 29.8000 ;
	    RECT 19.8000 28.8000 20.2000 29.2000 ;
         LAYER metal3 ;
	    RECT 19.8000 30.1500 20.2000 30.2000 ;
	    RECT 21.4000 30.1500 21.8000 30.2000 ;
	    RECT 19.8000 29.8500 21.8000 30.1500 ;
	    RECT 19.8000 29.8000 20.2000 29.8500 ;
	    RECT 21.4000 29.8000 21.8000 29.8500 ;
      END
   END s[6]
   PIN s[5]
      PORT
         LAYER metal1 ;
	    RECT 0.6000 6.2000 1.0000 9.9000 ;
	    RECT 0.6000 5.1000 0.9000 6.2000 ;
	    RECT 0.6000 1.1000 1.0000 5.1000 ;
         LAYER metal2 ;
	    RECT 0.6000 4.8000 1.0000 5.2000 ;
	    RECT 0.6500 4.2000 0.9500 4.8000 ;
	    RECT 0.6000 3.8000 1.0000 4.2000 ;
         LAYER metal3 ;
	    RECT 0.6000 5.1500 1.0000 5.2000 ;
	    RECT -2.5500 4.8500 1.0000 5.1500 ;
	    RECT 0.6000 4.8000 1.0000 4.8500 ;
      END
   END s[5]
   PIN s[4]
      PORT
         LAYER metal1 ;
	    RECT 0.6000 26.2000 1.0000 29.9000 ;
	    RECT 0.6000 25.1000 0.9000 26.2000 ;
	    RECT 0.6000 21.1000 1.0000 25.1000 ;
         LAYER metal2 ;
	    RECT 0.6000 24.8000 1.0000 25.2000 ;
	    RECT 0.6500 24.2000 0.9500 24.8000 ;
	    RECT 0.6000 23.8000 1.0000 24.2000 ;
         LAYER metal3 ;
	    RECT 0.6000 25.1500 1.0000 25.2000 ;
	    RECT -2.5500 24.8500 1.0000 25.1500 ;
	    RECT 0.6000 24.8000 1.0000 24.8500 ;
      END
   END s[4]
   PIN s[3]
      PORT
         LAYER metal1 ;
	    RECT 27.0000 6.2000 27.4000 9.9000 ;
	    RECT 27.0000 5.1000 27.3000 6.2000 ;
	    RECT 27.0000 1.1000 27.4000 5.1000 ;
         LAYER metal2 ;
	    RECT 27.0000 1.8000 27.4000 2.2000 ;
	    RECT 27.0500 -1.8500 27.3500 1.8000 ;
	    RECT 27.0500 -2.1500 28.1500 -1.8500 ;
      END
   END s[3]
   PIN s[2]
      PORT
         LAYER metal1 ;
	    RECT 60.6000 26.2000 61.0000 29.9000 ;
	    RECT 60.7000 25.1000 61.0000 26.2000 ;
	    RECT 60.6000 21.1000 61.0000 25.1000 ;
         LAYER metal2 ;
	    RECT 59.8500 33.8500 60.9500 34.1500 ;
	    RECT 60.6500 29.2000 60.9500 33.8500 ;
	    RECT 60.6000 28.8000 61.0000 29.2000 ;
      END
   END s[2]
   PIN s[1]
      PORT
         LAYER metal1 ;
	    RECT 63.8000 15.9000 64.2000 19.9000 ;
	    RECT 63.9000 14.8000 64.2000 15.9000 ;
	    RECT 63.8000 14.1500 64.2000 14.8000 ;
	    RECT 64.6000 14.1500 65.0000 14.2000 ;
	    RECT 63.8000 13.8500 65.0000 14.1500 ;
	    RECT 63.8000 11.1000 64.2000 13.8500 ;
	    RECT 64.6000 13.8000 65.0000 13.8500 ;
         LAYER metal2 ;
	    RECT 64.6000 14.8000 65.0000 15.2000 ;
	    RECT 64.6500 14.2000 64.9500 14.8000 ;
	    RECT 64.6000 13.8000 65.0000 14.2000 ;
         LAYER metal3 ;
	    RECT 64.6000 15.1500 65.0000 15.2000 ;
	    RECT 64.6000 14.8500 67.3500 15.1500 ;
	    RECT 64.6000 14.8000 65.0000 14.8500 ;
      END
   END s[1]
   PIN s[0]
      PORT
         LAYER metal1 ;
	    RECT 63.0000 26.2000 63.4000 29.9000 ;
	    RECT 63.1000 25.1000 63.4000 26.2000 ;
	    RECT 63.0000 24.1500 63.4000 25.1000 ;
	    RECT 64.6000 24.1500 65.0000 24.2000 ;
	    RECT 63.0000 23.8500 65.0000 24.1500 ;
	    RECT 63.0000 21.1000 63.4000 23.8500 ;
	    RECT 64.6000 23.8000 65.0000 23.8500 ;
         LAYER metal2 ;
	    RECT 64.6000 24.8000 65.0000 25.2000 ;
	    RECT 64.6500 24.2000 64.9500 24.8000 ;
	    RECT 64.6000 23.8000 65.0000 24.2000 ;
         LAYER metal3 ;
	    RECT 64.6000 25.1500 65.0000 25.2000 ;
	    RECT 64.6000 24.8500 67.3500 25.1500 ;
	    RECT 64.6000 24.8000 65.0000 24.8500 ;
      END
   END s[0]
   PIN x[5]
      PORT
         LAYER metal1 ;
	    RECT 0.6000 13.8000 1.4000 14.2000 ;
	    RECT 6.2000 12.4000 6.6000 13.2000 ;
         LAYER metal2 ;
	    RECT 0.6000 13.8000 1.0000 14.2000 ;
	    RECT 0.6500 13.2000 0.9500 13.8000 ;
	    RECT 0.6000 12.8000 1.0000 13.2000 ;
	    RECT 6.2000 13.1500 6.6000 13.2000 ;
	    RECT 7.0000 13.1500 7.4000 13.2000 ;
	    RECT 6.2000 12.8500 7.4000 13.1500 ;
	    RECT 6.2000 12.8000 6.6000 12.8500 ;
	    RECT 7.0000 12.8000 7.4000 12.8500 ;
         LAYER metal3 ;
	    RECT 0.6000 14.1500 1.0000 14.2000 ;
	    RECT -2.5500 13.8500 1.0000 14.1500 ;
	    RECT 0.6000 13.8000 1.0000 13.8500 ;
	    RECT 0.6000 13.1500 1.0000 13.2000 ;
	    RECT 7.0000 13.1500 7.4000 13.2000 ;
	    RECT 0.6000 12.8500 7.4000 13.1500 ;
	    RECT 0.6000 12.8000 1.0000 12.8500 ;
	    RECT 7.0000 12.8000 7.4000 12.8500 ;
      END
   END x[5]
   PIN x[4]
      PORT
         LAYER metal1 ;
	    RECT 14.2000 27.8000 14.6000 28.6000 ;
	    RECT 13.0000 27.1500 13.8000 27.2000 ;
	    RECT 14.2500 27.1500 14.5500 27.8000 ;
	    RECT 13.0000 26.8500 14.5500 27.1500 ;
	    RECT 13.0000 26.8000 13.8000 26.8500 ;
         LAYER metal2 ;
	    RECT 14.2500 28.2000 14.5500 34.1500 ;
	    RECT 14.2000 27.8000 14.6000 28.2000 ;
      END
   END x[4]
   PIN x[3]
      PORT
         LAYER metal1 ;
	    RECT 31.8000 27.8000 32.2000 28.6000 ;
	    RECT 26.6000 26.8000 27.4000 27.2000 ;
         LAYER metal2 ;
	    RECT 31.8500 28.2000 32.1500 34.1500 ;
	    RECT 27.0000 27.8000 27.4000 28.2000 ;
	    RECT 31.8000 27.8000 32.2000 28.2000 ;
	    RECT 27.0500 27.2000 27.3500 27.8000 ;
	    RECT 27.0000 26.8000 27.4000 27.2000 ;
         LAYER metal3 ;
	    RECT 27.0000 28.1500 27.4000 28.2000 ;
	    RECT 31.8000 28.1500 32.2000 28.2000 ;
	    RECT 27.0000 27.8500 32.2000 28.1500 ;
	    RECT 27.0000 27.8000 27.4000 27.8500 ;
	    RECT 31.8000 27.8000 32.2000 27.8500 ;
      END
   END x[3]
   PIN x[2]
      PORT
         LAYER metal1 ;
	    RECT 43.0000 27.8000 43.4000 28.6000 ;
	    RECT 43.0500 27.1500 43.3500 27.8000 ;
	    RECT 43.8000 27.1500 44.6000 27.2000 ;
	    RECT 43.0500 26.8500 44.6000 27.1500 ;
	    RECT 43.8000 26.8000 44.6000 26.8500 ;
         LAYER metal2 ;
	    RECT 43.8500 27.2000 44.1500 34.1500 ;
	    RECT 43.8000 26.8000 44.2000 27.2000 ;
      END
   END x[2]
   PIN x[1]
      PORT
         LAYER metal1 ;
	    RECT 44.6000 8.1500 45.0000 8.6000 ;
	    RECT 44.6000 7.8500 47.3500 8.1500 ;
	    RECT 44.6000 7.8000 45.0000 7.8500 ;
	    RECT 47.0500 7.1500 47.3500 7.8500 ;
	    RECT 47.8000 7.1500 48.6000 7.2000 ;
	    RECT 47.0500 6.8500 48.6000 7.1500 ;
	    RECT 47.8000 6.8000 48.6000 6.8500 ;
	    RECT 47.8500 6.1500 48.1500 6.8000 ;
	    RECT 49.4000 6.1500 49.8000 6.2000 ;
	    RECT 47.8500 5.8500 49.8000 6.1500 ;
	    RECT 49.4000 5.8000 49.8000 5.8500 ;
         LAYER metal2 ;
	    RECT 49.4000 5.8000 49.8000 6.2000 ;
	    RECT 49.4500 -2.1500 49.7500 5.8000 ;
      END
   END x[1]
   PIN x[0]
      PORT
         LAYER metal1 ;
	    RECT 58.2000 27.8000 58.6000 28.6000 ;
	    RECT 61.8000 7.1500 62.6000 7.2000 ;
	    RECT 63.0000 7.1500 63.4000 7.2000 ;
	    RECT 61.8000 6.8500 63.4000 7.1500 ;
	    RECT 61.8000 6.8000 62.6000 6.8500 ;
	    RECT 63.0000 6.8000 63.4000 6.8500 ;
         LAYER metal2 ;
	    RECT 58.2000 27.8000 58.6000 28.2000 ;
	    RECT 58.2500 27.1500 58.5500 27.8000 ;
	    RECT 58.2500 26.8500 59.3500 27.1500 ;
	    RECT 59.0500 18.2000 59.3500 26.8500 ;
	    RECT 59.0000 17.8000 59.4000 18.2000 ;
	    RECT 63.0000 17.8000 63.4000 18.2000 ;
	    RECT 63.0500 7.2000 63.3500 17.8000 ;
	    RECT 63.0000 6.8000 63.4000 7.2000 ;
         LAYER metal3 ;
	    RECT 59.0000 18.1500 59.4000 18.2000 ;
	    RECT 63.0000 18.1500 63.4000 18.2000 ;
	    RECT 59.0000 17.8500 67.3500 18.1500 ;
	    RECT 59.0000 17.8000 59.4000 17.8500 ;
	    RECT 63.0000 17.8000 63.4000 17.8500 ;
      END
   END x[0]
   PIN y[5]
      PORT
         LAYER metal1 ;
	    RECT 3.6000 14.3000 4.0000 14.4000 ;
	    RECT 3.6000 14.2000 5.0000 14.3000 ;
	    RECT 3.6000 14.0000 5.8000 14.2000 ;
	    RECT 4.7000 13.9000 5.8000 14.0000 ;
	    RECT 5.0000 13.8000 5.8000 13.9000 ;
	    RECT 7.8000 12.4000 8.2000 13.2000 ;
         LAYER metal2 ;
	    RECT 5.4000 15.8000 5.8000 16.2000 ;
	    RECT 5.4500 14.2000 5.7500 15.8000 ;
	    RECT 5.4000 14.1500 5.8000 14.2000 ;
	    RECT 6.2000 14.1500 6.6000 14.2000 ;
	    RECT 5.4000 13.8500 6.6000 14.1500 ;
	    RECT 5.4000 13.8000 5.8000 13.8500 ;
	    RECT 6.2000 13.8000 6.6000 13.8500 ;
	    RECT 7.8000 13.8000 8.2000 14.2000 ;
	    RECT 7.8500 13.2000 8.1500 13.8000 ;
	    RECT 7.8000 12.8000 8.2000 13.2000 ;
         LAYER metal3 ;
	    RECT 5.4000 16.1500 5.8000 16.2000 ;
	    RECT -2.5500 15.8500 5.8000 16.1500 ;
	    RECT 5.4000 15.8000 5.8000 15.8500 ;
	    RECT 6.2000 14.1500 6.6000 14.2000 ;
	    RECT 7.8000 14.1500 8.2000 14.2000 ;
	    RECT 6.2000 13.8500 8.2000 14.1500 ;
	    RECT 6.2000 13.8000 6.6000 13.8500 ;
	    RECT 7.8000 13.8000 8.2000 13.8500 ;
      END
   END y[5]
   PIN y[4]
      PORT
         LAYER metal1 ;
	    RECT 15.8000 27.8000 16.2000 28.6000 ;
	    RECT 8.6000 27.1000 9.4000 27.2000 ;
	    RECT 8.6000 27.0000 9.7000 27.1000 ;
	    RECT 8.6000 26.8000 10.8000 27.0000 ;
	    RECT 9.4000 26.7000 10.8000 26.8000 ;
	    RECT 10.4000 26.6000 10.8000 26.7000 ;
         LAYER metal2 ;
	    RECT 19.8500 31.2000 20.1500 34.1500 ;
	    RECT 8.6000 30.8000 9.0000 31.2000 ;
	    RECT 15.8000 30.8000 16.2000 31.2000 ;
	    RECT 19.8000 30.8000 20.2000 31.2000 ;
	    RECT 8.6500 27.2000 8.9500 30.8000 ;
	    RECT 15.8500 28.2000 16.1500 30.8000 ;
	    RECT 15.8000 27.8000 16.2000 28.2000 ;
	    RECT 8.6000 26.8000 9.0000 27.2000 ;
         LAYER metal3 ;
	    RECT 8.6000 31.1500 9.0000 31.2000 ;
	    RECT 15.8000 31.1500 16.2000 31.2000 ;
	    RECT 19.8000 31.1500 20.2000 31.2000 ;
	    RECT 8.6000 30.8500 20.2000 31.1500 ;
	    RECT 8.6000 30.8000 9.0000 30.8500 ;
	    RECT 15.8000 30.8000 16.2000 30.8500 ;
	    RECT 19.8000 30.8000 20.2000 30.8500 ;
      END
   END y[4]
   PIN y[3]
      PORT
         LAYER metal1 ;
	    RECT 27.8000 27.8000 28.2000 28.6000 ;
	    RECT 22.2000 27.1000 23.0000 27.2000 ;
	    RECT 22.2000 27.0000 23.3000 27.1000 ;
	    RECT 22.2000 26.8000 24.4000 27.0000 ;
	    RECT 23.0000 26.7000 24.4000 26.8000 ;
	    RECT 24.0000 26.6000 24.4000 26.7000 ;
         LAYER metal2 ;
	    RECT 27.8500 28.2000 28.1500 34.1500 ;
	    RECT 22.2000 27.8000 22.6000 28.2000 ;
	    RECT 27.8000 27.8000 28.2000 28.2000 ;
	    RECT 22.2500 27.2000 22.5500 27.8000 ;
	    RECT 27.8500 27.2000 28.1500 27.8000 ;
	    RECT 22.2000 26.8000 22.6000 27.2000 ;
	    RECT 27.8000 26.8000 28.2000 27.2000 ;
         LAYER metal3 ;
	    RECT 22.2000 27.8000 22.6000 28.2000 ;
	    RECT 22.2500 27.1500 22.5500 27.8000 ;
	    RECT 27.8000 27.1500 28.2000 27.2000 ;
	    RECT 22.2500 26.8500 28.2000 27.1500 ;
	    RECT 27.8000 26.8000 28.2000 26.8500 ;
      END
   END y[3]
   PIN y[2]
      PORT
         LAYER metal1 ;
	    RECT 41.4000 27.8000 41.8000 28.6000 ;
	    RECT 48.2000 27.1000 49.0000 27.2000 ;
	    RECT 47.9000 27.0000 49.0000 27.1000 ;
	    RECT 46.8000 26.8000 49.0000 27.0000 ;
	    RECT 46.8000 26.7000 48.2000 26.8000 ;
	    RECT 46.8000 26.6000 47.2000 26.7000 ;
         LAYER metal2 ;
	    RECT 41.4500 28.2000 41.7500 34.1500 ;
	    RECT 41.4000 27.8000 41.8000 28.2000 ;
	    RECT 48.6000 27.8000 49.0000 28.2000 ;
	    RECT 41.4500 27.2000 41.7500 27.8000 ;
	    RECT 48.6500 27.2000 48.9500 27.8000 ;
	    RECT 41.4000 26.8000 41.8000 27.2000 ;
	    RECT 48.6000 26.8000 49.0000 27.2000 ;
         LAYER metal3 ;
	    RECT 48.6000 27.8000 49.0000 28.2000 ;
	    RECT 41.4000 27.1500 41.8000 27.2000 ;
	    RECT 48.6500 27.1500 48.9500 27.8000 ;
	    RECT 41.4000 26.8500 48.9500 27.1500 ;
	    RECT 41.4000 26.8000 41.8000 26.8500 ;
      END
   END y[2]
   PIN y[1]
      PORT
         LAYER metal1 ;
	    RECT 38.2000 7.8000 38.6000 8.6000 ;
	    RECT 52.2000 7.1000 53.0000 7.2000 ;
	    RECT 51.9000 7.0000 53.0000 7.1000 ;
	    RECT 50.8000 6.8000 53.0000 7.0000 ;
	    RECT 50.8000 6.7000 52.2000 6.8000 ;
	    RECT 50.8000 6.6000 51.2000 6.7000 ;
         LAYER metal2 ;
	    RECT 38.2000 8.1500 38.6000 8.2000 ;
	    RECT 39.0000 8.1500 39.4000 8.2000 ;
	    RECT 38.2000 7.8500 39.4000 8.1500 ;
	    RECT 38.2000 7.8000 38.6000 7.8500 ;
	    RECT 39.0000 7.8000 39.4000 7.8500 ;
	    RECT 52.6000 7.8000 53.0000 8.2000 ;
	    RECT 52.6500 7.2000 52.9500 7.8000 ;
	    RECT 52.6000 6.8000 53.0000 7.2000 ;
	    RECT 52.6500 1.2000 52.9500 6.8000 ;
	    RECT 51.0000 0.8000 51.4000 1.2000 ;
	    RECT 52.6000 0.8000 53.0000 1.2000 ;
	    RECT 51.0500 -2.1500 51.3500 0.8000 ;
         LAYER metal3 ;
	    RECT 39.0000 8.1500 39.4000 8.2000 ;
	    RECT 52.6000 8.1500 53.0000 8.2000 ;
	    RECT 38.2500 7.8500 53.0000 8.1500 ;
	    RECT 39.0000 7.8000 39.4000 7.8500 ;
	    RECT 52.6000 7.8000 53.0000 7.8500 ;
	    RECT 51.0000 1.1500 51.4000 1.2000 ;
	    RECT 52.6000 1.1500 53.0000 1.2000 ;
	    RECT 51.0000 0.8500 53.0000 1.1500 ;
	    RECT 51.0000 0.8000 51.4000 0.8500 ;
	    RECT 52.6000 0.8000 53.0000 0.8500 ;
      END
   END y[1]
   PIN y[0]
      PORT
         LAYER metal1 ;
	    RECT 54.2000 7.8000 54.6000 8.6000 ;
	    RECT 57.4000 7.1000 58.2000 7.2000 ;
	    RECT 57.4000 7.0000 58.5000 7.1000 ;
	    RECT 57.4000 6.8000 59.6000 7.0000 ;
	    RECT 58.2000 6.7000 59.6000 6.8000 ;
	    RECT 59.2000 6.6000 59.6000 6.7000 ;
         LAYER metal2 ;
	    RECT 54.2000 7.8000 54.6000 8.2000 ;
	    RECT 54.2500 7.2000 54.5500 7.8000 ;
	    RECT 54.2000 6.8000 54.6000 7.2000 ;
	    RECT 56.6000 7.1500 57.0000 7.2000 ;
	    RECT 57.4000 7.1500 57.8000 7.2000 ;
	    RECT 56.6000 6.8500 57.8000 7.1500 ;
	    RECT 56.6000 6.8000 57.0000 6.8500 ;
	    RECT 57.4000 6.8000 57.8000 6.8500 ;
	    RECT 57.4500 1.2000 57.7500 6.8000 ;
	    RECT 57.4000 0.8000 57.8000 1.2000 ;
	    RECT 59.0000 0.8000 59.4000 1.2000 ;
	    RECT 59.0500 -2.1500 59.3500 0.8000 ;
         LAYER metal3 ;
	    RECT 54.2000 7.1500 54.6000 7.2000 ;
	    RECT 56.6000 7.1500 57.0000 7.2000 ;
	    RECT 54.2000 6.8500 57.0000 7.1500 ;
	    RECT 54.2000 6.8000 54.6000 6.8500 ;
	    RECT 56.6000 6.8000 57.0000 6.8500 ;
	    RECT 57.4000 1.1500 57.8000 1.2000 ;
	    RECT 59.0000 1.1500 59.4000 1.2000 ;
	    RECT 57.4000 0.8500 59.4000 1.1500 ;
	    RECT 57.4000 0.8000 57.8000 0.8500 ;
	    RECT 59.0000 0.8000 59.4000 0.8500 ;
      END
   END y[0]
   OBS
         LAYER metal1 ;
	    RECT 2.2000 27.6000 2.6000 29.9000 ;
	    RECT 3.0000 27.9000 3.4000 29.9000 ;
	    RECT 5.2000 28.1000 6.0000 29.9000 ;
	    RECT 3.0000 27.6000 4.3000 27.9000 ;
	    RECT 1.5000 27.3000 2.6000 27.6000 ;
	    RECT 3.9000 27.5000 4.3000 27.6000 ;
	    RECT 4.6000 27.4000 5.4000 27.8000 ;
	    RECT 1.5000 25.8000 1.8000 27.3000 ;
	    RECT 3.0000 27.1000 3.8000 27.2000 ;
	    RECT 5.7000 27.1000 6.0000 28.1000 ;
	    RECT 7.8000 27.9000 8.2000 29.9000 ;
	    RECT 6.3000 27.4000 6.7000 27.8000 ;
	    RECT 7.0000 27.6000 8.2000 27.9000 ;
	    RECT 8.6000 27.9000 9.0000 29.9000 ;
	    RECT 10.8000 29.2000 11.6000 29.9000 ;
	    RECT 10.2000 28.8000 11.6000 29.2000 ;
	    RECT 10.8000 28.1000 11.6000 28.8000 ;
	    RECT 8.6000 27.6000 9.9000 27.9000 ;
	    RECT 7.0000 27.5000 7.4000 27.6000 ;
	    RECT 9.5000 27.5000 9.9000 27.6000 ;
	    RECT 10.2000 27.4000 11.0000 27.8000 ;
	    RECT 3.0000 27.0000 4.1000 27.1000 ;
	    RECT 3.0000 26.8000 5.2000 27.0000 ;
	    RECT 3.8000 26.7000 5.2000 26.8000 ;
	    RECT 4.8000 26.6000 5.2000 26.7000 ;
	    RECT 5.5000 26.8000 6.0000 27.1000 ;
	    RECT 6.4000 27.2000 6.7000 27.4000 ;
	    RECT 6.4000 26.8000 6.8000 27.2000 ;
	    RECT 7.4000 26.8000 8.2000 27.2000 ;
	    RECT 11.3000 27.1000 11.6000 28.1000 ;
	    RECT 13.4000 27.9000 13.8000 29.9000 ;
	    RECT 11.9000 27.4000 12.3000 27.8000 ;
	    RECT 12.6000 27.6000 13.8000 27.9000 ;
	    RECT 12.6000 27.5000 13.0000 27.6000 ;
	    RECT 11.1000 26.8000 11.6000 27.1000 ;
	    RECT 12.0000 27.2000 12.3000 27.4000 ;
	    RECT 12.0000 26.8000 12.4000 27.2000 ;
	    RECT 2.2000 25.8000 2.6000 26.6000 ;
	    RECT 5.5000 26.2000 5.8000 26.8000 ;
	    RECT 11.1000 26.2000 11.4000 26.8000 ;
	    RECT 4.1000 26.1000 4.5000 26.2000 ;
	    RECT 4.1000 25.8000 4.9000 26.1000 ;
	    RECT 5.4000 25.8000 5.8000 26.2000 ;
	    RECT 9.7000 26.1000 10.1000 26.2000 ;
	    RECT 9.7000 25.8000 10.5000 26.1000 ;
	    RECT 11.0000 25.8000 11.4000 26.2000 ;
	    RECT 1.2000 25.4000 1.8000 25.8000 ;
	    RECT 4.5000 25.7000 4.9000 25.8000 ;
	    RECT 1.5000 25.1000 1.8000 25.4000 ;
	    RECT 5.5000 25.1000 5.8000 25.8000 ;
	    RECT 10.1000 25.7000 10.5000 25.8000 ;
	    RECT 11.1000 25.1000 11.4000 25.8000 ;
	    RECT 1.5000 24.8000 2.6000 25.1000 ;
	    RECT 2.2000 21.1000 2.6000 24.8000 ;
	    RECT 3.0000 24.8000 4.3000 25.1000 ;
	    RECT 3.0000 21.1000 3.4000 24.8000 ;
	    RECT 3.9000 24.7000 4.3000 24.8000 ;
	    RECT 5.2000 21.1000 6.0000 25.1000 ;
	    RECT 7.0000 24.8000 8.2000 25.1000 ;
	    RECT 7.0000 24.7000 7.4000 24.8000 ;
	    RECT 7.8000 21.1000 8.2000 24.8000 ;
	    RECT 8.6000 24.8000 9.9000 25.1000 ;
	    RECT 8.6000 21.1000 9.0000 24.8000 ;
	    RECT 9.5000 24.7000 9.9000 24.8000 ;
	    RECT 10.8000 21.1000 11.6000 25.1000 ;
	    RECT 12.6000 24.8000 13.8000 25.1000 ;
	    RECT 12.6000 24.7000 13.0000 24.8000 ;
	    RECT 13.4000 21.1000 13.8000 24.8000 ;
	    RECT 14.2000 24.1500 14.6000 24.2000 ;
	    RECT 15.0000 24.1500 15.4000 29.9000 ;
	    RECT 14.2000 23.8500 15.4000 24.1500 ;
	    RECT 14.2000 23.8000 14.6000 23.8500 ;
	    RECT 15.0000 21.1000 15.4000 23.8500 ;
	    RECT 16.6000 22.1500 17.0000 29.9000 ;
	    RECT 21.4000 27.6000 21.8000 29.9000 ;
	    RECT 22.2000 27.9000 22.6000 29.9000 ;
	    RECT 24.4000 28.1000 25.2000 29.9000 ;
	    RECT 22.2000 27.6000 23.5000 27.9000 ;
	    RECT 20.7000 27.3000 21.8000 27.6000 ;
	    RECT 23.1000 27.5000 23.5000 27.6000 ;
	    RECT 23.8000 27.4000 24.6000 27.8000 ;
	    RECT 20.7000 25.8000 21.0000 27.3000 ;
	    RECT 24.9000 27.1000 25.2000 28.1000 ;
	    RECT 27.0000 27.9000 27.4000 29.9000 ;
	    RECT 25.5000 27.4000 25.9000 27.8000 ;
	    RECT 26.2000 27.6000 27.4000 27.9000 ;
	    RECT 28.6000 28.1500 29.0000 29.9000 ;
	    RECT 30.2000 28.9000 30.6000 29.9000 ;
	    RECT 29.4000 28.1500 29.8000 28.6000 ;
	    RECT 28.6000 27.8500 29.8000 28.1500 ;
	    RECT 26.2000 27.5000 26.6000 27.6000 ;
	    RECT 24.7000 26.8000 25.2000 27.1000 ;
	    RECT 25.6000 27.2000 25.9000 27.4000 ;
	    RECT 25.6000 26.8000 26.0000 27.2000 ;
	    RECT 28.6000 27.1500 29.0000 27.8500 ;
	    RECT 29.4000 27.8000 29.8000 27.8500 ;
	    RECT 30.3000 27.2000 30.6000 28.9000 ;
	    RECT 28.6000 26.8500 29.7500 27.1500 ;
	    RECT 21.4000 25.8000 21.8000 26.6000 ;
	    RECT 24.7000 26.2000 25.0000 26.8000 ;
	    RECT 23.3000 26.1000 23.7000 26.2000 ;
	    RECT 23.3000 25.8000 24.1000 26.1000 ;
	    RECT 24.6000 25.8000 25.0000 26.2000 ;
	    RECT 20.4000 25.4000 21.0000 25.8000 ;
	    RECT 23.7000 25.7000 24.1000 25.8000 ;
	    RECT 20.7000 25.1000 21.0000 25.4000 ;
	    RECT 24.7000 25.1000 25.0000 25.8000 ;
	    RECT 20.7000 24.8000 21.8000 25.1000 ;
	    RECT 18.2000 22.1500 18.6000 22.2000 ;
	    RECT 16.6000 21.8500 18.6000 22.1500 ;
	    RECT 16.6000 21.1000 17.0000 21.8500 ;
	    RECT 18.2000 21.8000 18.6000 21.8500 ;
	    RECT 21.4000 21.1000 21.8000 24.8000 ;
	    RECT 22.2000 24.8000 23.5000 25.1000 ;
	    RECT 22.2000 21.1000 22.6000 24.8000 ;
	    RECT 23.1000 24.7000 23.5000 24.8000 ;
	    RECT 24.4000 22.2000 25.2000 25.1000 ;
	    RECT 26.2000 24.8000 27.4000 25.1000 ;
	    RECT 26.2000 24.7000 26.6000 24.8000 ;
	    RECT 24.4000 21.8000 25.8000 22.2000 ;
	    RECT 24.4000 21.1000 25.2000 21.8000 ;
	    RECT 27.0000 21.1000 27.4000 24.8000 ;
	    RECT 28.6000 21.1000 29.0000 26.8500 ;
	    RECT 29.4500 26.2000 29.7500 26.8500 ;
	    RECT 30.2000 26.8000 30.6000 27.2000 ;
	    RECT 29.4000 25.8000 29.8000 26.2000 ;
	    RECT 30.3000 25.1000 30.6000 26.8000 ;
	    RECT 31.0000 26.1500 31.4000 26.2000 ;
	    RECT 32.6000 26.1500 33.0000 29.9000 ;
	    RECT 33.7000 28.2000 34.1000 29.9000 ;
	    RECT 36.6000 28.9000 37.0000 29.9000 ;
	    RECT 33.7000 27.9000 34.6000 28.2000 ;
	    RECT 31.0000 25.8500 33.0000 26.1500 ;
	    RECT 31.0000 25.4000 31.4000 25.8500 ;
	    RECT 32.6000 25.1500 33.0000 25.8500 ;
	    RECT 33.4000 26.1500 33.8000 26.2000 ;
	    RECT 34.2000 26.1500 34.6000 27.9000 ;
	    RECT 35.0000 26.8000 35.4000 27.6000 ;
	    RECT 36.6000 27.2000 36.9000 28.9000 ;
	    RECT 37.4000 27.8000 37.8000 28.6000 ;
	    RECT 38.5000 28.2000 38.9000 29.9000 ;
	    RECT 38.5000 27.9000 39.4000 28.2000 ;
	    RECT 36.6000 26.8000 37.0000 27.2000 ;
	    RECT 33.4000 25.8500 34.6000 26.1500 ;
	    RECT 33.4000 25.8000 33.8000 25.8500 ;
	    RECT 33.4000 25.1500 33.8000 25.2000 ;
	    RECT 30.2000 24.7000 31.1000 25.1000 ;
	    RECT 30.7000 22.2000 31.1000 24.7000 ;
	    RECT 30.2000 21.8000 31.1000 22.2000 ;
	    RECT 30.7000 21.1000 31.1000 21.8000 ;
	    RECT 32.6000 24.8500 33.8000 25.1500 ;
	    RECT 32.6000 21.1000 33.0000 24.8500 ;
	    RECT 33.4000 24.4000 33.8000 24.8500 ;
	    RECT 34.2000 21.1000 34.6000 25.8500 ;
	    RECT 35.8000 25.4000 36.2000 26.2000 ;
	    RECT 36.6000 25.1000 36.9000 26.8000 ;
	    RECT 36.1000 24.7000 37.0000 25.1000 ;
	    RECT 36.1000 22.2000 36.5000 24.7000 ;
	    RECT 38.2000 24.4000 38.6000 25.2000 ;
	    RECT 35.8000 21.8000 36.5000 22.2000 ;
	    RECT 36.1000 21.1000 36.5000 21.8000 ;
	    RECT 39.0000 24.1500 39.4000 27.9000 ;
	    RECT 39.8000 27.1500 40.2000 27.6000 ;
	    RECT 40.6000 27.1500 41.0000 29.9000 ;
	    RECT 39.8000 26.8500 41.0000 27.1500 ;
	    RECT 39.8000 26.8000 40.2000 26.8500 ;
	    RECT 39.8000 24.1500 40.2000 24.2000 ;
	    RECT 39.0000 23.8500 40.2000 24.1500 ;
	    RECT 39.0000 21.1000 39.4000 23.8500 ;
	    RECT 39.8000 23.8000 40.2000 23.8500 ;
	    RECT 40.6000 21.1000 41.0000 26.8500 ;
	    RECT 41.4000 25.8000 41.8000 26.2000 ;
	    RECT 41.4500 25.1500 41.7500 25.8000 ;
	    RECT 42.2000 25.1500 42.6000 29.9000 ;
	    RECT 43.8000 27.9000 44.2000 29.9000 ;
	    RECT 46.0000 28.1000 46.8000 29.9000 ;
	    RECT 43.8000 27.6000 45.0000 27.9000 ;
	    RECT 44.6000 27.5000 45.0000 27.6000 ;
	    RECT 45.3000 27.4000 45.7000 27.8000 ;
	    RECT 45.3000 27.2000 45.6000 27.4000 ;
	    RECT 45.2000 26.8000 45.6000 27.2000 ;
	    RECT 46.0000 27.1000 46.3000 28.1000 ;
	    RECT 48.6000 27.9000 49.0000 29.9000 ;
	    RECT 46.6000 27.4000 47.4000 27.8000 ;
	    RECT 47.7000 27.6000 49.0000 27.9000 ;
	    RECT 51.8000 27.9000 52.2000 29.9000 ;
	    RECT 54.0000 28.1000 54.8000 29.9000 ;
	    RECT 51.8000 27.6000 53.0000 27.9000 ;
	    RECT 47.7000 27.5000 48.1000 27.6000 ;
	    RECT 52.6000 27.5000 53.0000 27.6000 ;
	    RECT 53.3000 27.4000 53.7000 27.8000 ;
	    RECT 53.3000 27.2000 53.6000 27.4000 ;
	    RECT 46.0000 26.8000 46.5000 27.1000 ;
	    RECT 51.8000 26.8000 52.6000 27.2000 ;
	    RECT 53.2000 26.8000 53.6000 27.2000 ;
	    RECT 54.0000 27.1000 54.3000 28.1000 ;
	    RECT 56.6000 27.9000 57.0000 29.9000 ;
	    RECT 54.6000 27.4000 55.4000 27.8000 ;
	    RECT 55.7000 27.6000 57.0000 27.9000 ;
	    RECT 55.7000 27.5000 56.1000 27.6000 ;
	    RECT 56.2000 27.1000 57.0000 27.2000 ;
	    RECT 54.0000 26.8000 54.5000 27.1000 ;
	    RECT 55.9000 27.0000 57.0000 27.1000 ;
	    RECT 46.2000 26.2000 46.5000 26.8000 ;
	    RECT 54.2000 26.2000 54.5000 26.8000 ;
	    RECT 54.8000 26.8000 57.0000 27.0000 ;
	    RECT 54.8000 26.7000 56.2000 26.8000 ;
	    RECT 54.8000 26.6000 55.2000 26.7000 ;
	    RECT 45.4000 26.1500 45.8000 26.2000 ;
	    RECT 46.2000 26.1500 46.6000 26.2000 ;
	    RECT 45.4000 25.8500 46.6000 26.1500 ;
	    RECT 47.5000 26.1000 47.9000 26.2000 ;
	    RECT 45.4000 25.8000 45.8000 25.8500 ;
	    RECT 46.2000 25.8000 46.6000 25.8500 ;
	    RECT 47.1000 25.8000 47.9000 26.1000 ;
	    RECT 54.2000 25.8000 54.6000 26.2000 ;
	    RECT 55.5000 26.1000 55.9000 26.2000 ;
	    RECT 55.1000 25.8000 55.9000 26.1000 ;
	    RECT 41.4500 24.8500 42.6000 25.1500 ;
	    RECT 46.2000 25.1000 46.5000 25.8000 ;
	    RECT 47.1000 25.7000 47.5000 25.8000 ;
	    RECT 54.2000 25.1000 54.5000 25.8000 ;
	    RECT 55.1000 25.7000 55.5000 25.8000 ;
	    RECT 42.2000 21.1000 42.6000 24.8500 ;
	    RECT 43.8000 24.8000 45.0000 25.1000 ;
	    RECT 43.8000 21.1000 44.2000 24.8000 ;
	    RECT 44.6000 24.7000 45.0000 24.8000 ;
	    RECT 46.0000 21.1000 46.8000 25.1000 ;
	    RECT 47.7000 24.8000 49.0000 25.1000 ;
	    RECT 47.7000 24.7000 48.1000 24.8000 ;
	    RECT 48.6000 21.1000 49.0000 24.8000 ;
	    RECT 51.8000 24.8000 53.0000 25.1000 ;
	    RECT 51.8000 21.1000 52.2000 24.8000 ;
	    RECT 52.6000 24.7000 53.0000 24.8000 ;
	    RECT 54.0000 21.1000 54.8000 25.1000 ;
	    RECT 55.7000 24.8000 57.0000 25.1000 ;
	    RECT 55.7000 24.7000 56.1000 24.8000 ;
	    RECT 56.6000 21.1000 57.0000 24.8000 ;
	    RECT 57.4000 21.1000 57.8000 29.9000 ;
	    RECT 59.0000 27.6000 59.4000 29.9000 ;
	    RECT 61.4000 27.6000 61.8000 29.9000 ;
	    RECT 59.0000 27.3000 60.1000 27.6000 ;
	    RECT 61.4000 27.3000 62.5000 27.6000 ;
	    RECT 59.0000 26.1500 59.4000 26.6000 ;
	    RECT 58.2500 25.8500 59.4000 26.1500 ;
	    RECT 58.2500 25.2000 58.5500 25.8500 ;
	    RECT 59.0000 25.8000 59.4000 25.8500 ;
	    RECT 59.8000 25.8000 60.1000 27.3000 ;
	    RECT 61.4000 25.8000 61.8000 26.6000 ;
	    RECT 62.2000 25.8000 62.5000 27.3000 ;
	    RECT 59.8000 25.4000 60.4000 25.8000 ;
	    RECT 62.2000 25.4000 62.8000 25.8000 ;
	    RECT 58.2000 24.8000 58.6000 25.2000 ;
	    RECT 59.8000 25.1000 60.1000 25.4000 ;
	    RECT 62.2000 25.1000 62.5000 25.4000 ;
	    RECT 59.0000 24.8000 60.1000 25.1000 ;
	    RECT 61.4000 24.8000 62.5000 25.1000 ;
	    RECT 59.0000 21.1000 59.4000 24.8000 ;
	    RECT 61.4000 21.1000 61.8000 24.8000 ;
	    RECT 0.6000 16.2000 1.0000 19.9000 ;
	    RECT 1.4000 16.2000 1.8000 16.3000 ;
	    RECT 0.6000 15.9000 1.8000 16.2000 ;
	    RECT 2.8000 15.9000 3.6000 19.9000 ;
	    RECT 4.5000 16.2000 4.9000 16.3000 ;
	    RECT 5.4000 16.2000 5.8000 19.9000 ;
	    RECT 4.5000 15.9000 5.8000 16.2000 ;
	    RECT 3.0000 15.2000 3.3000 15.9000 ;
	    RECT 3.9000 15.2000 4.3000 15.3000 ;
	    RECT 3.0000 14.8000 3.4000 15.2000 ;
	    RECT 3.9000 14.9000 4.7000 15.2000 ;
	    RECT 4.3000 14.8000 4.7000 14.9000 ;
	    RECT 7.0000 15.1500 7.4000 19.9000 ;
	    RECT 7.8000 15.8000 8.2000 16.2000 ;
	    RECT 7.8500 15.1500 8.1500 15.8000 ;
	    RECT 7.0000 14.8500 8.1500 15.1500 ;
	    RECT 3.0000 14.2000 3.3000 14.8000 ;
	    RECT 2.0000 13.8000 2.4000 14.2000 ;
	    RECT 2.1000 13.6000 2.4000 13.8000 ;
	    RECT 2.8000 13.9000 3.3000 14.2000 ;
	    RECT 1.4000 13.4000 1.8000 13.5000 ;
	    RECT 0.6000 13.1000 1.8000 13.4000 ;
	    RECT 2.1000 13.2000 2.5000 13.6000 ;
	    RECT 0.6000 11.1000 1.0000 13.1000 ;
	    RECT 2.8000 12.9000 3.1000 13.9000 ;
	    RECT 3.4000 13.2000 4.2000 13.6000 ;
	    RECT 4.5000 13.4000 4.9000 13.5000 ;
	    RECT 4.5000 13.1000 5.8000 13.4000 ;
	    RECT 2.8000 11.1000 3.6000 12.9000 ;
	    RECT 5.4000 11.1000 5.8000 13.1000 ;
	    RECT 7.0000 11.1000 7.4000 14.8500 ;
	    RECT 8.6000 13.1500 9.0000 19.9000 ;
	    RECT 9.7000 16.3000 10.1000 19.9000 ;
	    RECT 9.7000 15.9000 10.6000 16.3000 ;
	    RECT 9.4000 14.8000 9.8000 15.6000 ;
	    RECT 10.2000 14.2000 10.5000 15.9000 ;
	    RECT 9.4000 13.8000 9.8000 14.2000 ;
	    RECT 10.2000 13.8000 10.6000 14.2000 ;
	    RECT 11.8000 14.1500 12.2000 14.2000 ;
	    RECT 11.0500 13.8500 12.2000 14.1500 ;
	    RECT 9.4500 13.1500 9.7500 13.8000 ;
	    RECT 8.6000 12.8500 9.7500 13.1500 ;
	    RECT 8.6000 11.1000 9.0000 12.8500 ;
	    RECT 10.2000 12.2000 10.5000 13.8000 ;
	    RECT 11.0500 13.2000 11.3500 13.8500 ;
	    RECT 11.8000 13.4000 12.2000 13.8500 ;
	    RECT 11.0000 12.4000 11.4000 13.2000 ;
	    RECT 12.6000 13.1000 13.0000 19.9000 ;
	    RECT 13.4000 15.8000 13.8000 16.6000 ;
	    RECT 14.2000 15.8000 14.6000 16.6000 ;
	    RECT 15.0000 13.1000 15.4000 19.9000 ;
	    RECT 19.3000 16.3000 19.7000 19.9000 ;
	    RECT 19.3000 15.9000 20.2000 16.3000 ;
	    RECT 19.0000 14.8000 19.4000 15.6000 ;
	    RECT 19.8000 14.2000 20.1000 15.9000 ;
	    RECT 15.8000 13.4000 16.2000 14.2000 ;
	    RECT 19.8000 14.1500 20.2000 14.2000 ;
	    RECT 21.4000 14.1500 21.8000 14.2000 ;
	    RECT 19.8000 13.8500 21.8000 14.1500 ;
	    RECT 19.8000 13.8000 20.2000 13.8500 ;
	    RECT 12.6000 12.8000 13.5000 13.1000 ;
	    RECT 13.1000 12.2000 13.5000 12.8000 ;
	    RECT 14.5000 12.8000 15.4000 13.1000 ;
	    RECT 14.5000 12.2000 14.9000 12.8000 ;
	    RECT 19.8000 12.2000 20.1000 13.8000 ;
	    RECT 21.4000 13.4000 21.8000 13.8500 ;
	    RECT 20.6000 12.4000 21.0000 13.2000 ;
	    RECT 22.2000 13.1000 22.6000 19.9000 ;
	    RECT 23.0000 15.8000 23.4000 16.6000 ;
	    RECT 24.6000 14.1500 25.0000 19.9000 ;
	    RECT 25.4000 14.1500 25.8000 14.2000 ;
	    RECT 24.6000 13.8500 25.8000 14.1500 ;
	    RECT 22.2000 12.8000 23.1000 13.1000 ;
	    RECT 10.2000 11.1000 10.6000 12.2000 ;
	    RECT 13.1000 11.8000 13.8000 12.2000 ;
	    RECT 14.5000 11.8000 15.4000 12.2000 ;
	    RECT 13.1000 11.1000 13.5000 11.8000 ;
	    RECT 14.5000 11.1000 14.9000 11.8000 ;
	    RECT 19.8000 11.1000 20.2000 12.2000 ;
	    RECT 22.7000 11.1000 23.1000 12.8000 ;
	    RECT 23.8000 12.4000 24.2000 13.2000 ;
	    RECT 24.6000 11.1000 25.0000 13.8500 ;
	    RECT 25.4000 13.4000 25.8000 13.8500 ;
	    RECT 26.2000 13.1000 26.6000 19.9000 ;
	    RECT 27.0000 15.8000 27.4000 16.6000 ;
	    RECT 27.8000 16.2000 28.2000 19.9000 ;
	    RECT 28.6000 16.2000 29.0000 16.3000 ;
	    RECT 27.8000 15.9000 29.0000 16.2000 ;
	    RECT 30.0000 15.9000 30.8000 19.9000 ;
	    RECT 31.7000 16.2000 32.1000 16.3000 ;
	    RECT 32.6000 16.2000 33.0000 19.9000 ;
	    RECT 31.7000 15.9000 33.0000 16.2000 ;
	    RECT 30.2000 15.2000 30.5000 15.9000 ;
	    RECT 33.4000 15.8000 33.8000 16.6000 ;
	    RECT 31.1000 15.2000 31.5000 15.3000 ;
	    RECT 30.2000 14.8000 30.6000 15.2000 ;
	    RECT 31.1000 14.9000 31.9000 15.2000 ;
	    RECT 31.5000 14.8000 31.9000 14.9000 ;
	    RECT 30.2000 14.2000 30.5000 14.8000 ;
	    RECT 27.8000 13.8000 28.6000 14.2000 ;
	    RECT 29.2000 13.8000 29.6000 14.2000 ;
	    RECT 29.3000 13.6000 29.6000 13.8000 ;
	    RECT 30.0000 13.9000 30.5000 14.2000 ;
	    RECT 30.8000 14.3000 31.2000 14.4000 ;
	    RECT 30.8000 14.2000 32.2000 14.3000 ;
	    RECT 30.8000 14.0000 33.0000 14.2000 ;
	    RECT 31.9000 13.9000 33.0000 14.0000 ;
	    RECT 28.6000 13.4000 29.0000 13.5000 ;
	    RECT 27.8000 13.1000 29.0000 13.4000 ;
	    RECT 29.3000 13.2000 29.7000 13.6000 ;
	    RECT 26.2000 12.8000 27.1000 13.1000 ;
	    RECT 26.7000 12.2000 27.1000 12.8000 ;
	    RECT 26.2000 11.8000 27.1000 12.2000 ;
	    RECT 26.7000 11.1000 27.1000 11.8000 ;
	    RECT 27.8000 11.1000 28.2000 13.1000 ;
	    RECT 30.0000 12.9000 30.3000 13.9000 ;
	    RECT 32.2000 13.8000 33.0000 13.9000 ;
	    RECT 30.6000 13.2000 31.4000 13.6000 ;
	    RECT 31.7000 13.4000 32.1000 13.5000 ;
	    RECT 31.7000 13.1000 33.0000 13.4000 ;
	    RECT 34.2000 13.1000 34.6000 19.9000 ;
	    RECT 35.0000 14.1500 35.4000 14.2000 ;
	    RECT 35.8000 14.1500 36.2000 14.2000 ;
	    RECT 35.0000 13.8500 36.2000 14.1500 ;
	    RECT 35.0000 13.4000 35.4000 13.8500 ;
	    RECT 35.8000 13.8000 36.2000 13.8500 ;
	    RECT 36.6000 14.1500 37.0000 19.9000 ;
	    RECT 37.4000 14.1500 37.8000 14.2000 ;
	    RECT 36.6000 13.8500 37.8000 14.1500 ;
	    RECT 30.0000 11.1000 30.8000 12.9000 ;
	    RECT 32.6000 11.1000 33.0000 13.1000 ;
	    RECT 33.7000 12.8000 34.6000 13.1000 ;
	    RECT 33.7000 12.2000 34.1000 12.8000 ;
	    RECT 35.8000 12.4000 36.2000 13.2000 ;
	    RECT 33.4000 11.8000 34.1000 12.2000 ;
	    RECT 33.7000 11.1000 34.1000 11.8000 ;
	    RECT 36.6000 11.1000 37.0000 13.8500 ;
	    RECT 37.4000 13.4000 37.8000 13.8500 ;
	    RECT 38.2000 13.1000 38.6000 19.9000 ;
	    RECT 40.6000 17.9000 41.0000 19.9000 ;
	    RECT 39.0000 15.8000 39.4000 16.6000 ;
	    RECT 40.7000 15.8000 41.0000 17.9000 ;
	    RECT 42.2000 15.9000 42.6000 19.9000 ;
	    RECT 40.7000 15.5000 41.9000 15.8000 ;
	    RECT 40.6000 14.8000 41.0000 15.2000 ;
	    RECT 39.8000 13.8000 40.2000 14.6000 ;
	    RECT 40.7000 14.4000 41.0000 14.8000 ;
	    RECT 40.7000 14.1000 41.2000 14.4000 ;
	    RECT 40.8000 14.0000 41.2000 14.1000 ;
	    RECT 41.6000 13.8000 41.9000 15.5000 ;
	    RECT 42.3000 15.2000 42.6000 15.9000 ;
	    RECT 43.0000 15.8000 43.4000 16.6000 ;
	    RECT 42.2000 14.8000 42.6000 15.2000 ;
	    RECT 43.8000 15.1500 44.2000 19.9000 ;
	    RECT 45.4000 15.8000 45.8000 16.6000 ;
	    RECT 41.6000 13.7000 42.0000 13.8000 ;
	    RECT 40.5000 13.5000 42.0000 13.7000 ;
	    RECT 39.9000 13.4000 42.0000 13.5000 ;
	    RECT 39.9000 13.2000 40.8000 13.4000 ;
	    RECT 39.9000 13.1000 40.2000 13.2000 ;
	    RECT 42.3000 13.1000 42.6000 14.8000 ;
	    RECT 43.0500 14.8500 44.2000 15.1500 ;
	    RECT 43.0500 14.2000 43.3500 14.8500 ;
	    RECT 43.0000 13.8000 43.4000 14.2000 ;
	    RECT 43.8000 13.1000 44.2000 14.8500 ;
	    RECT 44.6000 13.4000 45.0000 14.2000 ;
	    RECT 46.2000 13.1000 46.6000 19.9000 ;
	    RECT 47.0000 13.4000 47.4000 14.2000 ;
	    RECT 51.0000 14.1500 51.4000 19.9000 ;
	    RECT 51.8000 14.1500 52.2000 14.2000 ;
	    RECT 51.0000 13.8500 52.2000 14.1500 ;
	    RECT 38.2000 12.8000 39.1000 13.1000 ;
	    RECT 38.7000 11.1000 39.1000 12.8000 ;
	    RECT 39.8000 11.1000 40.2000 13.1000 ;
	    RECT 41.9000 12.6000 42.6000 13.1000 ;
	    RECT 43.3000 12.8000 44.2000 13.1000 ;
	    RECT 45.7000 12.8000 46.6000 13.1000 ;
	    RECT 41.9000 11.1000 42.3000 12.6000 ;
	    RECT 43.3000 11.1000 43.7000 12.8000 ;
	    RECT 45.7000 12.2000 46.1000 12.8000 ;
	    RECT 50.2000 12.4000 50.6000 13.2000 ;
	    RECT 45.4000 11.8000 46.1000 12.2000 ;
	    RECT 45.7000 11.1000 46.1000 11.8000 ;
	    RECT 51.0000 11.1000 51.4000 13.8500 ;
	    RECT 51.8000 13.4000 52.2000 13.8500 ;
	    RECT 52.6000 14.1500 53.0000 19.9000 ;
	    RECT 53.4000 15.8000 53.8000 16.6000 ;
	    RECT 54.2000 15.8000 54.6000 16.6000 ;
	    RECT 53.4500 15.1500 53.7500 15.8000 ;
	    RECT 55.0000 15.1500 55.4000 19.9000 ;
	    RECT 56.6000 16.2000 57.0000 19.9000 ;
	    RECT 57.4000 16.2000 57.8000 16.3000 ;
	    RECT 56.6000 15.9000 57.8000 16.2000 ;
	    RECT 58.8000 15.9000 59.6000 19.9000 ;
	    RECT 60.5000 16.2000 60.9000 16.3000 ;
	    RECT 61.4000 16.2000 61.8000 19.9000 ;
	    RECT 60.5000 15.9000 61.8000 16.2000 ;
	    RECT 62.2000 16.2000 62.6000 19.9000 ;
	    RECT 62.2000 15.9000 63.3000 16.2000 ;
	    RECT 53.4500 14.8500 55.4000 15.1500 ;
	    RECT 53.4000 14.1500 53.8000 14.2000 ;
	    RECT 52.6000 13.8500 53.8000 14.1500 ;
	    RECT 52.6000 13.1000 53.0000 13.8500 ;
	    RECT 53.4000 13.8000 53.8000 13.8500 ;
	    RECT 55.0000 13.1000 55.4000 14.8500 ;
	    RECT 59.0000 15.8000 59.4000 15.9000 ;
	    RECT 59.0000 15.2000 59.3000 15.8000 ;
	    RECT 63.0000 15.6000 63.3000 15.9000 ;
	    RECT 59.9000 15.2000 60.3000 15.3000 ;
	    RECT 63.0000 15.2000 63.6000 15.6000 ;
	    RECT 59.0000 14.8000 59.4000 15.2000 ;
	    RECT 59.9000 14.9000 60.7000 15.2000 ;
	    RECT 60.3000 14.8000 60.7000 14.9000 ;
	    RECT 59.0000 14.2000 59.3000 14.8000 ;
	    RECT 62.2000 14.4000 62.6000 15.2000 ;
	    RECT 55.8000 13.4000 56.2000 14.2000 ;
	    RECT 56.6000 13.8000 57.4000 14.2000 ;
	    RECT 58.0000 13.8000 58.4000 14.2000 ;
	    RECT 58.1000 13.6000 58.4000 13.8000 ;
	    RECT 58.8000 13.9000 59.3000 14.2000 ;
	    RECT 59.6000 14.3000 60.0000 14.4000 ;
	    RECT 59.6000 14.2000 61.0000 14.3000 ;
	    RECT 59.6000 14.0000 61.8000 14.2000 ;
	    RECT 60.7000 13.9000 61.8000 14.0000 ;
	    RECT 57.4000 13.4000 57.8000 13.5000 ;
	    RECT 52.6000 12.8000 53.5000 13.1000 ;
	    RECT 53.1000 11.1000 53.5000 12.8000 ;
	    RECT 54.5000 12.8000 55.4000 13.1000 ;
	    RECT 56.6000 13.1000 57.8000 13.4000 ;
	    RECT 58.1000 13.2000 58.5000 13.6000 ;
	    RECT 54.5000 11.1000 54.9000 12.8000 ;
	    RECT 56.6000 11.1000 57.0000 13.1000 ;
	    RECT 58.8000 12.9000 59.1000 13.9000 ;
	    RECT 61.0000 13.8000 61.8000 13.9000 ;
	    RECT 63.0000 13.7000 63.3000 15.2000 ;
	    RECT 59.4000 13.2000 60.2000 13.6000 ;
	    RECT 60.5000 13.4000 60.9000 13.5000 ;
	    RECT 62.2000 13.4000 63.3000 13.7000 ;
	    RECT 60.5000 13.1000 61.8000 13.4000 ;
	    RECT 58.8000 11.1000 59.6000 12.9000 ;
	    RECT 61.4000 11.1000 61.8000 13.1000 ;
	    RECT 62.2000 11.1000 62.6000 13.4000 ;
	    RECT 2.2000 7.6000 2.6000 9.9000 ;
	    RECT 3.0000 7.9000 3.4000 9.9000 ;
	    RECT 5.2000 8.1000 6.0000 9.9000 ;
	    RECT 3.0000 7.6000 4.2000 7.9000 ;
	    RECT 1.5000 7.3000 2.6000 7.6000 ;
	    RECT 3.8000 7.5000 4.2000 7.6000 ;
	    RECT 4.5000 7.4000 4.9000 7.8000 ;
	    RECT 1.5000 5.8000 1.8000 7.3000 ;
	    RECT 4.5000 7.2000 4.8000 7.4000 ;
	    RECT 3.0000 6.8000 3.8000 7.2000 ;
	    RECT 4.4000 6.8000 4.8000 7.2000 ;
	    RECT 5.2000 7.1000 5.5000 8.1000 ;
	    RECT 7.8000 7.9000 8.2000 9.9000 ;
	    RECT 9.9000 8.2000 10.3000 9.9000 ;
	    RECT 5.8000 7.4000 6.6000 7.8000 ;
	    RECT 6.9000 7.6000 8.2000 7.9000 ;
	    RECT 9.4000 7.9000 10.3000 8.2000 ;
	    RECT 11.3000 8.2000 11.7000 9.9000 ;
	    RECT 11.3000 7.9000 12.2000 8.2000 ;
	    RECT 6.9000 7.5000 7.3000 7.6000 ;
	    RECT 7.4000 7.1000 8.2000 7.2000 ;
	    RECT 5.2000 6.8000 5.7000 7.1000 ;
	    RECT 7.1000 7.0000 8.2000 7.1000 ;
	    RECT 2.2000 6.1500 2.6000 6.6000 ;
	    RECT 5.4000 6.2000 5.7000 6.8000 ;
	    RECT 6.0000 6.8000 8.2000 7.0000 ;
	    RECT 8.6000 6.8000 9.0000 7.6000 ;
	    RECT 6.0000 6.7000 7.4000 6.8000 ;
	    RECT 6.0000 6.6000 6.4000 6.7000 ;
	    RECT 5.4000 6.1500 5.8000 6.2000 ;
	    RECT 2.2000 5.8500 5.8000 6.1500 ;
	    RECT 6.7000 6.1000 7.1000 6.2000 ;
	    RECT 2.2000 5.8000 2.6000 5.8500 ;
	    RECT 5.4000 5.8000 5.8000 5.8500 ;
	    RECT 6.3000 5.8000 7.1000 6.1000 ;
	    RECT 9.4000 6.1500 9.8000 7.9000 ;
	    RECT 11.0000 7.1500 11.4000 7.2000 ;
	    RECT 11.8000 7.1500 12.2000 7.9000 ;
	    RECT 11.0000 6.8500 12.2000 7.1500 ;
	    RECT 11.0000 6.8000 11.4000 6.8500 ;
	    RECT 9.4000 5.8500 11.3500 6.1500 ;
	    RECT 1.2000 5.4000 1.8000 5.8000 ;
	    RECT 1.5000 5.1000 1.8000 5.4000 ;
	    RECT 5.4000 5.1000 5.7000 5.8000 ;
	    RECT 6.3000 5.7000 6.7000 5.8000 ;
	    RECT 1.5000 4.8000 2.6000 5.1000 ;
	    RECT 2.2000 1.1000 2.6000 4.8000 ;
	    RECT 3.0000 4.8000 4.2000 5.1000 ;
	    RECT 3.0000 1.1000 3.4000 4.8000 ;
	    RECT 3.8000 4.7000 4.2000 4.8000 ;
	    RECT 5.2000 1.1000 6.0000 5.1000 ;
	    RECT 6.9000 4.8000 8.2000 5.1000 ;
	    RECT 6.9000 4.7000 7.3000 4.8000 ;
	    RECT 7.8000 1.1000 8.2000 4.8000 ;
	    RECT 9.4000 1.1000 9.8000 5.8500 ;
	    RECT 11.0500 5.2000 11.3500 5.8500 ;
	    RECT 10.2000 4.4000 10.6000 5.2000 ;
	    RECT 11.0000 4.4000 11.4000 5.2000 ;
	    RECT 11.8000 1.1000 12.2000 6.8500 ;
	    RECT 12.6000 7.1500 13.0000 7.6000 ;
	    RECT 13.4000 7.1500 13.8000 9.9000 ;
	    RECT 14.2000 7.8000 14.6000 8.6000 ;
	    RECT 15.0000 7.9000 15.4000 9.9000 ;
	    RECT 17.1000 8.4000 17.5000 9.9000 ;
	    RECT 17.1000 7.9000 17.8000 8.4000 ;
	    RECT 20.9000 8.2000 21.3000 9.9000 ;
	    RECT 23.3000 9.2000 23.7000 9.9000 ;
	    RECT 23.0000 8.8000 23.7000 9.2000 ;
	    RECT 23.3000 8.2000 23.7000 8.8000 ;
	    RECT 20.9000 7.9000 21.8000 8.2000 ;
	    RECT 23.3000 7.9000 24.2000 8.2000 ;
	    RECT 15.1000 7.8000 15.4000 7.9000 ;
	    RECT 15.1000 7.6000 16.0000 7.8000 ;
	    RECT 15.1000 7.5000 17.2000 7.6000 ;
	    RECT 15.7000 7.3000 17.2000 7.5000 ;
	    RECT 16.8000 7.2000 17.2000 7.3000 ;
	    RECT 12.6000 6.8500 13.8000 7.1500 ;
	    RECT 12.6000 6.8000 13.0000 6.8500 ;
	    RECT 13.4000 1.1000 13.8000 6.8500 ;
	    RECT 14.2000 7.1500 14.6000 7.2000 ;
	    RECT 15.0000 7.1500 15.4000 7.2000 ;
	    RECT 14.2000 6.8500 15.4000 7.1500 ;
	    RECT 16.0000 6.9000 16.4000 7.0000 ;
	    RECT 14.2000 6.8000 14.6000 6.8500 ;
	    RECT 15.0000 6.4000 15.4000 6.8500 ;
	    RECT 15.9000 6.6000 16.4000 6.9000 ;
	    RECT 15.9000 6.2000 16.2000 6.6000 ;
	    RECT 15.8000 5.8000 16.2000 6.2000 ;
	    RECT 16.8000 5.5000 17.1000 7.2000 ;
	    RECT 17.5000 6.2000 17.8000 7.9000 ;
	    RECT 17.4000 5.8000 17.8000 6.2000 ;
	    RECT 15.9000 5.2000 17.1000 5.5000 ;
	    RECT 15.9000 3.1000 16.2000 5.2000 ;
	    RECT 17.5000 5.1500 17.8000 5.8000 ;
	    RECT 20.6000 5.1500 21.0000 5.2000 ;
	    RECT 17.4500 5.1000 21.0000 5.1500 ;
	    RECT 15.8000 1.1000 16.2000 3.1000 ;
	    RECT 17.4000 4.8500 21.0000 5.1000 ;
	    RECT 17.4000 1.1000 17.8000 4.8500 ;
	    RECT 20.6000 4.4000 21.0000 4.8500 ;
	    RECT 21.4000 5.1500 21.8000 7.9000 ;
	    RECT 22.2000 6.8000 22.6000 7.6000 ;
	    RECT 23.0000 5.1500 23.4000 5.2000 ;
	    RECT 21.4000 4.8500 23.4000 5.1500 ;
	    RECT 21.4000 1.1000 21.8000 4.8500 ;
	    RECT 23.0000 4.4000 23.4000 4.8500 ;
	    RECT 23.8000 1.1000 24.2000 7.9000 ;
	    RECT 24.6000 7.1500 25.0000 7.6000 ;
	    RECT 25.4000 7.1500 25.8000 9.9000 ;
	    RECT 26.2000 7.8000 26.6000 8.6000 ;
	    RECT 28.6000 7.6000 29.0000 9.9000 ;
	    RECT 29.4000 7.8000 29.8000 8.6000 ;
	    RECT 24.6000 6.8500 25.8000 7.1500 ;
	    RECT 24.6000 6.8000 25.0000 6.8500 ;
	    RECT 25.4000 1.1000 25.8000 6.8500 ;
	    RECT 27.9000 7.3000 29.0000 7.6000 ;
	    RECT 27.9000 5.8000 28.2000 7.3000 ;
	    RECT 30.2000 7.1500 30.6000 9.9000 ;
	    RECT 32.3000 8.2000 32.7000 9.9000 ;
	    RECT 31.8000 8.1500 32.7000 8.2000 ;
	    RECT 33.4000 8.1500 33.8000 8.6000 ;
	    RECT 31.8000 7.8500 33.8000 8.1500 ;
	    RECT 31.0000 7.1500 31.4000 7.6000 ;
	    RECT 30.2000 6.8500 31.4000 7.1500 ;
	    RECT 28.6000 6.1500 29.0000 6.6000 ;
	    RECT 29.4000 6.1500 29.8000 6.2000 ;
	    RECT 28.6000 5.8500 29.8000 6.1500 ;
	    RECT 28.6000 5.8000 29.0000 5.8500 ;
	    RECT 29.4000 5.8000 29.8000 5.8500 ;
	    RECT 27.6000 5.4000 28.2000 5.8000 ;
	    RECT 27.9000 5.1000 28.2000 5.4000 ;
	    RECT 27.9000 4.8000 29.0000 5.1000 ;
	    RECT 28.6000 1.1000 29.0000 4.8000 ;
	    RECT 30.2000 1.1000 30.6000 6.8500 ;
	    RECT 31.0000 6.8000 31.4000 6.8500 ;
	    RECT 31.8000 1.1000 32.2000 7.8500 ;
	    RECT 33.4000 7.8000 33.8000 7.8500 ;
	    RECT 34.2000 7.1500 34.6000 9.9000 ;
	    RECT 36.3000 8.2000 36.7000 9.9000 ;
	    RECT 35.8000 7.9000 36.7000 8.2000 ;
	    RECT 35.0000 7.1500 35.4000 7.6000 ;
	    RECT 34.2000 6.8500 35.4000 7.1500 ;
	    RECT 32.6000 5.1500 33.0000 5.2000 ;
	    RECT 33.4000 5.1500 33.8000 5.2000 ;
	    RECT 32.6000 4.8500 33.8000 5.1500 ;
	    RECT 32.6000 4.4000 33.0000 4.8500 ;
	    RECT 33.4000 4.8000 33.8000 4.8500 ;
	    RECT 34.2000 1.1000 34.6000 6.8500 ;
	    RECT 35.0000 6.8000 35.4000 6.8500 ;
	    RECT 35.8000 1.1000 36.2000 7.9000 ;
	    RECT 37.4000 7.1500 37.8000 9.9000 ;
	    RECT 39.8000 8.8000 40.2000 9.9000 ;
	    RECT 39.0000 7.8000 39.4000 8.6000 ;
	    RECT 39.0500 7.1500 39.3500 7.8000 ;
	    RECT 39.9000 7.2000 40.2000 8.8000 ;
	    RECT 42.7000 9.2000 43.1000 9.9000 ;
	    RECT 42.7000 8.8000 43.4000 9.2000 ;
	    RECT 42.7000 8.2000 43.1000 8.8000 ;
	    RECT 42.2000 7.9000 43.1000 8.2000 ;
	    RECT 37.4000 6.8500 39.3500 7.1500 ;
	    RECT 36.6000 4.4000 37.0000 5.2000 ;
	    RECT 37.4000 1.1000 37.8000 6.8500 ;
	    RECT 39.0500 6.2000 39.3500 6.8500 ;
	    RECT 39.8000 6.8000 40.2000 7.2000 ;
	    RECT 41.4000 6.8000 41.8000 7.6000 ;
	    RECT 39.0000 5.8000 39.4000 6.2000 ;
	    RECT 39.9000 5.1000 40.2000 6.8000 ;
	    RECT 40.6000 5.4000 41.0000 6.2000 ;
	    RECT 39.8000 4.7000 40.7000 5.1000 ;
	    RECT 40.3000 1.1000 40.7000 4.7000 ;
	    RECT 42.2000 1.1000 42.6000 7.9000 ;
	    RECT 43.0000 6.8000 43.4000 7.2000 ;
	    RECT 43.0500 6.1500 43.3500 6.8000 ;
	    RECT 43.8000 6.1500 44.2000 9.9000 ;
	    RECT 47.8000 7.9000 48.2000 9.9000 ;
	    RECT 50.0000 9.2000 50.8000 9.9000 ;
	    RECT 50.0000 8.8000 51.4000 9.2000 ;
	    RECT 50.0000 8.1000 50.8000 8.8000 ;
	    RECT 47.8000 7.6000 49.0000 7.9000 ;
	    RECT 48.6000 7.5000 49.0000 7.6000 ;
	    RECT 49.3000 7.4000 49.7000 7.8000 ;
	    RECT 49.3000 7.2000 49.6000 7.4000 ;
	    RECT 49.2000 6.8000 49.6000 7.2000 ;
	    RECT 50.0000 7.1000 50.3000 8.1000 ;
	    RECT 52.6000 7.9000 53.0000 9.9000 ;
	    RECT 50.6000 7.4000 51.4000 7.8000 ;
	    RECT 51.7000 7.6000 53.0000 7.9000 ;
	    RECT 51.7000 7.5000 52.1000 7.6000 ;
	    RECT 53.4000 7.1500 53.8000 9.9000 ;
	    RECT 55.8000 8.8000 56.2000 9.9000 ;
	    RECT 55.0000 7.8000 55.4000 8.6000 ;
	    RECT 55.0500 7.1500 55.3500 7.8000 ;
	    RECT 55.9000 7.2000 56.2000 8.8000 ;
	    RECT 57.4000 7.9000 57.8000 9.9000 ;
	    RECT 59.6000 8.1000 60.4000 9.9000 ;
	    RECT 57.4000 7.6000 58.7000 7.9000 ;
	    RECT 58.3000 7.5000 58.7000 7.6000 ;
	    RECT 59.0000 7.4000 59.8000 7.8000 ;
	    RECT 50.0000 6.8000 50.5000 7.1000 ;
	    RECT 43.0500 5.8500 44.2000 6.1500 ;
	    RECT 43.0000 5.1500 43.4000 5.2000 ;
	    RECT 43.8000 5.1500 44.2000 5.8500 ;
	    RECT 43.0000 4.8500 44.2000 5.1500 ;
	    RECT 50.2000 6.2000 50.5000 6.8000 ;
	    RECT 53.4000 6.8500 55.3500 7.1500 ;
	    RECT 50.2000 5.8000 50.6000 6.2000 ;
	    RECT 51.5000 6.1000 51.9000 6.2000 ;
	    RECT 51.1000 5.8000 51.9000 6.1000 ;
	    RECT 50.2000 5.1000 50.5000 5.8000 ;
	    RECT 51.1000 5.7000 51.5000 5.8000 ;
	    RECT 43.0000 4.4000 43.4000 4.8500 ;
	    RECT 43.8000 1.1000 44.2000 4.8500 ;
	    RECT 47.8000 4.8000 49.0000 5.1000 ;
	    RECT 47.8000 1.1000 48.2000 4.8000 ;
	    RECT 48.6000 4.7000 49.0000 4.8000 ;
	    RECT 50.0000 1.1000 50.8000 5.1000 ;
	    RECT 51.7000 4.8000 53.0000 5.1000 ;
	    RECT 51.7000 4.7000 52.1000 4.8000 ;
	    RECT 52.6000 1.1000 53.0000 4.8000 ;
	    RECT 53.4000 1.1000 53.8000 6.8500 ;
	    RECT 55.8000 6.8000 56.2000 7.2000 ;
	    RECT 60.1000 7.1000 60.4000 8.1000 ;
	    RECT 62.2000 7.9000 62.6000 9.9000 ;
	    RECT 60.7000 7.4000 61.1000 7.8000 ;
	    RECT 61.4000 7.6000 62.6000 7.9000 ;
	    RECT 61.4000 7.5000 61.8000 7.6000 ;
	    RECT 55.9000 5.1000 56.2000 6.8000 ;
	    RECT 59.9000 6.8000 60.4000 7.1000 ;
	    RECT 60.8000 7.2000 61.1000 7.4000 ;
	    RECT 60.8000 6.8000 61.2000 7.2000 ;
	    RECT 59.9000 6.2000 60.2000 6.8000 ;
	    RECT 56.6000 5.4000 57.0000 6.2000 ;
	    RECT 58.5000 6.1000 58.9000 6.2000 ;
	    RECT 58.5000 5.8000 59.3000 6.1000 ;
	    RECT 59.8000 5.8000 60.2000 6.2000 ;
	    RECT 58.9000 5.7000 59.3000 5.8000 ;
	    RECT 59.9000 5.1000 60.2000 5.8000 ;
	    RECT 55.8000 4.7000 56.7000 5.1000 ;
	    RECT 56.3000 1.1000 56.7000 4.7000 ;
	    RECT 57.4000 4.8000 58.7000 5.1000 ;
	    RECT 57.4000 1.1000 57.8000 4.8000 ;
	    RECT 58.3000 4.7000 58.7000 4.8000 ;
	    RECT 59.6000 1.1000 60.4000 5.1000 ;
	    RECT 61.4000 4.8000 62.6000 5.1000 ;
	    RECT 61.4000 4.7000 61.8000 4.8000 ;
	    RECT 62.2000 1.1000 62.6000 4.8000 ;
         LAYER metal2 ;
	    RECT 7.8000 28.8000 8.2000 29.2000 ;
	    RECT 10.2000 29.1500 10.6000 29.2000 ;
	    RECT 11.0000 29.1500 11.4000 29.2000 ;
	    RECT 10.2000 28.8500 11.4000 29.1500 ;
	    RECT 10.2000 28.8000 10.6000 28.8500 ;
	    RECT 11.0000 28.8000 11.4000 28.8500 ;
	    RECT 3.9000 27.8000 4.3000 27.9000 ;
	    RECT 3.9000 27.5000 6.7000 27.8000 ;
	    RECT 7.0000 27.5000 7.4000 27.9000 ;
	    RECT 3.0000 26.8000 3.4000 27.2000 ;
	    RECT 1.4000 26.1500 1.8000 26.2000 ;
	    RECT 2.2000 26.1500 2.6000 26.2000 ;
	    RECT 1.4000 25.8500 2.6000 26.1500 ;
	    RECT 1.4000 25.8000 1.8000 25.8500 ;
	    RECT 2.2000 25.8000 2.6000 25.8500 ;
	    RECT 3.0500 25.2000 3.3500 26.8000 ;
	    RECT 3.0000 24.8000 3.4000 25.2000 ;
	    RECT 3.9000 25.1000 4.2000 27.5000 ;
	    RECT 4.6000 27.4000 5.0000 27.5000 ;
	    RECT 6.3000 27.4000 6.7000 27.5000 ;
	    RECT 7.1000 27.1000 7.4000 27.5000 ;
	    RECT 7.8500 27.2000 8.1500 28.8000 ;
	    RECT 37.4000 28.1500 37.8000 28.2000 ;
	    RECT 38.2000 28.1500 38.6000 28.2000 ;
	    RECT 9.5000 27.8000 9.9000 27.9000 ;
	    RECT 9.5000 27.5000 12.3000 27.8000 ;
	    RECT 12.6000 27.5000 13.0000 27.9000 ;
	    RECT 4.6000 26.8000 7.4000 27.1000 ;
	    RECT 7.8000 26.8000 8.2000 27.2000 ;
	    RECT 4.6000 26.1000 4.9000 26.8000 ;
	    RECT 4.5000 25.7000 4.9000 26.1000 ;
	    RECT 5.4000 25.8000 5.8000 26.2000 ;
	    RECT 5.4500 25.2000 5.7500 25.8000 ;
	    RECT 3.9000 24.7000 4.3000 25.1000 ;
	    RECT 5.4000 24.8000 5.8000 25.2000 ;
	    RECT 7.1000 25.1000 7.4000 26.8000 ;
	    RECT 7.0000 24.7000 7.4000 25.1000 ;
	    RECT 9.5000 25.1000 9.8000 27.5000 ;
	    RECT 10.2000 27.4000 10.6000 27.5000 ;
	    RECT 11.9000 27.4000 12.3000 27.5000 ;
	    RECT 12.7000 27.1000 13.0000 27.5000 ;
	    RECT 10.2000 26.8000 13.0000 27.1000 ;
	    RECT 10.2000 26.1000 10.5000 26.8000 ;
	    RECT 10.1000 25.7000 10.5000 26.1000 ;
	    RECT 12.7000 25.1000 13.0000 26.8000 ;
	    RECT 23.1000 27.8000 23.5000 27.9000 ;
	    RECT 23.1000 27.5000 25.9000 27.8000 ;
	    RECT 26.2000 27.5000 26.6000 27.9000 ;
	    RECT 37.4000 27.8500 38.6000 28.1500 ;
	    RECT 37.4000 27.8000 37.8000 27.8500 ;
	    RECT 38.2000 27.8000 38.6000 27.8500 ;
	    RECT 39.8000 27.8000 40.2000 28.2000 ;
	    RECT 21.4000 25.8000 21.8000 26.2000 ;
	    RECT 9.5000 24.7000 9.9000 25.1000 ;
	    RECT 12.6000 24.7000 13.0000 25.1000 ;
	    RECT 14.2000 23.8000 14.6000 24.2000 ;
	    RECT 1.4000 15.9000 1.8000 16.3000 ;
	    RECT 4.5000 15.9000 4.9000 16.3000 ;
	    RECT 14.2500 16.2000 14.5500 23.8000 ;
	    RECT 18.2000 22.1500 18.6000 22.2000 ;
	    RECT 19.0000 22.1500 19.4000 22.2000 ;
	    RECT 18.2000 21.8500 19.4000 22.1500 ;
	    RECT 18.2000 21.8000 18.6000 21.8500 ;
	    RECT 19.0000 21.8000 19.4000 21.8500 ;
	    RECT 20.6000 21.8000 21.0000 22.2000 ;
	    RECT 1.4000 14.2000 1.7000 15.9000 ;
	    RECT 3.9000 14.9000 4.3000 15.3000 ;
	    RECT 3.9000 14.2000 4.2000 14.9000 ;
	    RECT 1.4000 13.9000 4.2000 14.2000 ;
	    RECT 1.4000 13.5000 1.7000 13.9000 ;
	    RECT 2.1000 13.5000 2.5000 13.6000 ;
	    RECT 3.8000 13.5000 4.2000 13.6000 ;
	    RECT 4.6000 13.5000 4.9000 15.9000 ;
	    RECT 7.8000 15.8000 8.2000 16.2000 ;
	    RECT 13.4000 15.8000 13.8000 16.2000 ;
	    RECT 14.2000 15.8000 14.6000 16.2000 ;
	    RECT 7.8500 15.2000 8.1500 15.8000 ;
	    RECT 13.4500 15.2000 13.7500 15.8000 ;
	    RECT 14.2500 15.2000 14.5500 15.8000 ;
	    RECT 7.8000 14.8000 8.2000 15.2000 ;
	    RECT 8.6000 15.1500 9.0000 15.2000 ;
	    RECT 9.4000 15.1500 9.8000 15.2000 ;
	    RECT 8.6000 14.8500 9.8000 15.1500 ;
	    RECT 8.6000 14.8000 9.0000 14.8500 ;
	    RECT 9.4000 14.8000 9.8000 14.8500 ;
	    RECT 13.4000 14.8000 13.8000 15.2000 ;
	    RECT 14.2000 14.8000 14.6000 15.2000 ;
	    RECT 18.2000 15.1500 18.6000 15.2000 ;
	    RECT 19.0000 15.1500 19.4000 15.2000 ;
	    RECT 18.2000 14.8500 19.4000 15.1500 ;
	    RECT 18.2000 14.8000 18.6000 14.8500 ;
	    RECT 19.0000 14.8000 19.4000 14.8500 ;
	    RECT 20.6500 14.2000 20.9500 21.8000 ;
	    RECT 9.4000 13.8000 9.8000 14.2000 ;
	    RECT 15.8000 14.1500 16.2000 14.2000 ;
	    RECT 16.6000 14.1500 17.0000 14.2000 ;
	    RECT 15.8000 13.8500 17.0000 14.1500 ;
	    RECT 15.8000 13.8000 16.2000 13.8500 ;
	    RECT 16.6000 13.8000 17.0000 13.8500 ;
	    RECT 20.6000 13.8000 21.0000 14.2000 ;
	    RECT 1.4000 13.1000 1.8000 13.5000 ;
	    RECT 2.1000 13.2000 4.9000 13.5000 ;
	    RECT 9.4500 13.2000 9.7500 13.8000 ;
	    RECT 20.6500 13.2000 20.9500 13.8000 ;
	    RECT 4.5000 13.1000 4.9000 13.2000 ;
	    RECT 9.4000 12.8000 9.8000 13.2000 ;
	    RECT 10.2000 13.1500 10.6000 13.2000 ;
	    RECT 11.0000 13.1500 11.4000 13.2000 ;
	    RECT 10.2000 12.8500 11.4000 13.1500 ;
	    RECT 10.2000 12.8000 10.6000 12.8500 ;
	    RECT 11.0000 12.8000 11.4000 12.8500 ;
	    RECT 13.4000 12.8000 13.8000 13.2000 ;
	    RECT 20.6000 12.8000 21.0000 13.2000 ;
	    RECT 13.4500 12.2000 13.7500 12.8000 ;
	    RECT 3.0000 11.8000 3.4000 12.2000 ;
	    RECT 10.2000 12.1500 10.6000 12.2000 ;
	    RECT 11.0000 12.1500 11.4000 12.2000 ;
	    RECT 10.2000 11.8500 11.4000 12.1500 ;
	    RECT 10.2000 11.8000 10.6000 11.8500 ;
	    RECT 11.0000 11.8000 11.4000 11.8500 ;
	    RECT 13.4000 11.8000 13.8000 12.2000 ;
	    RECT 15.0000 11.8000 15.4000 12.2000 ;
	    RECT 19.8000 11.8000 20.2000 12.2000 ;
	    RECT 3.0500 7.2000 3.3500 11.8000 ;
	    RECT 3.8000 7.5000 4.2000 7.9000 ;
	    RECT 6.9000 7.8000 7.3000 7.9000 ;
	    RECT 8.6000 7.8000 9.0000 8.2000 ;
	    RECT 4.5000 7.5000 7.3000 7.8000 ;
	    RECT 3.0000 6.8000 3.4000 7.2000 ;
	    RECT 3.8000 7.1000 4.1000 7.5000 ;
	    RECT 4.5000 7.4000 4.9000 7.5000 ;
	    RECT 6.2000 7.4000 6.6000 7.5000 ;
	    RECT 3.8000 6.8000 6.6000 7.1000 ;
	    RECT 3.8000 5.1000 4.1000 6.8000 ;
	    RECT 6.3000 6.1000 6.6000 6.8000 ;
	    RECT 6.3000 5.7000 6.7000 6.1000 ;
	    RECT 7.0000 5.1000 7.3000 7.5000 ;
	    RECT 8.6500 7.2000 8.9500 7.8000 ;
	    RECT 7.8000 6.8000 8.2000 7.2000 ;
	    RECT 8.6000 6.8000 9.0000 7.2000 ;
	    RECT 10.2000 7.1500 10.6000 7.2000 ;
	    RECT 11.0000 7.1500 11.4000 7.2000 ;
	    RECT 10.2000 6.8500 11.4000 7.1500 ;
	    RECT 13.4500 7.1500 13.7500 11.8000 ;
	    RECT 14.2000 8.8000 14.6000 9.2000 ;
	    RECT 14.2500 8.2000 14.5500 8.8000 ;
	    RECT 14.2000 7.8000 14.6000 8.2000 ;
	    RECT 14.2000 7.1500 14.6000 7.2000 ;
	    RECT 13.4500 6.8500 14.6000 7.1500 ;
	    RECT 10.2000 6.8000 10.6000 6.8500 ;
	    RECT 11.0000 6.8000 11.4000 6.8500 ;
	    RECT 14.2000 6.8000 14.6000 6.8500 ;
	    RECT 7.8500 6.2000 8.1500 6.8000 ;
	    RECT 7.8000 5.8000 8.2000 6.2000 ;
	    RECT 15.0500 6.1500 15.3500 11.8000 ;
	    RECT 19.8500 9.2000 20.1500 11.8000 ;
	    RECT 21.4500 9.2000 21.7500 25.8000 ;
	    RECT 23.1000 25.1000 23.4000 27.5000 ;
	    RECT 23.8000 27.4000 24.2000 27.5000 ;
	    RECT 25.5000 27.4000 25.9000 27.5000 ;
	    RECT 26.3000 27.1000 26.6000 27.5000 ;
	    RECT 39.8500 27.2000 40.1500 27.8000 ;
	    RECT 44.6000 27.5000 45.0000 27.9000 ;
	    RECT 47.7000 27.8000 48.1000 27.9000 ;
	    RECT 45.3000 27.5000 48.1000 27.8000 ;
	    RECT 23.8000 26.8000 26.6000 27.1000 ;
	    RECT 29.4000 26.8000 29.8000 27.2000 ;
	    RECT 34.2000 27.1500 34.6000 27.2000 ;
	    RECT 35.0000 27.1500 35.4000 27.2000 ;
	    RECT 34.2000 26.8500 35.4000 27.1500 ;
	    RECT 34.2000 26.8000 34.6000 26.8500 ;
	    RECT 35.0000 26.8000 35.4000 26.8500 ;
	    RECT 39.8000 26.8000 40.2000 27.2000 ;
	    RECT 44.6000 27.1000 44.9000 27.5000 ;
	    RECT 45.3000 27.4000 45.7000 27.5000 ;
	    RECT 47.0000 27.4000 47.4000 27.5000 ;
	    RECT 44.6000 26.8000 47.4000 27.1000 ;
	    RECT 23.8000 26.1000 24.1000 26.8000 ;
	    RECT 23.7000 25.7000 24.1000 26.1000 ;
	    RECT 26.3000 25.1000 26.6000 26.8000 ;
	    RECT 29.4500 26.2000 29.7500 26.8000 ;
	    RECT 29.4000 25.8000 29.8000 26.2000 ;
	    RECT 33.4000 25.8000 33.8000 26.2000 ;
	    RECT 35.8000 25.8000 36.2000 26.2000 ;
	    RECT 41.4000 25.8000 41.8000 26.2000 ;
	    RECT 23.1000 24.7000 23.5000 25.1000 ;
	    RECT 26.2000 24.7000 26.6000 25.1000 ;
	    RECT 24.6000 22.1500 25.0000 22.2000 ;
	    RECT 25.4000 22.1500 25.8000 22.2000 ;
	    RECT 24.6000 21.8500 25.8000 22.1500 ;
	    RECT 24.6000 21.8000 25.0000 21.8500 ;
	    RECT 25.4000 21.8000 25.8000 21.8500 ;
	    RECT 27.8000 21.8000 28.2000 22.2000 ;
	    RECT 30.2000 21.8000 30.6000 22.2000 ;
	    RECT 22.2000 16.8000 22.6000 17.2000 ;
	    RECT 22.2500 16.2000 22.5500 16.8000 ;
	    RECT 22.2000 15.8000 22.6000 16.2000 ;
	    RECT 23.0000 15.8000 23.4000 16.2000 ;
	    RECT 26.2000 16.1500 26.6000 16.2000 ;
	    RECT 27.0000 16.1500 27.4000 16.2000 ;
	    RECT 26.2000 15.8500 27.4000 16.1500 ;
	    RECT 26.2000 15.8000 26.6000 15.8500 ;
	    RECT 27.0000 15.8000 27.4000 15.8500 ;
	    RECT 23.0500 13.2000 23.3500 15.8000 ;
	    RECT 27.8500 14.2000 28.1500 21.8000 ;
	    RECT 28.6000 15.9000 29.0000 16.3000 ;
	    RECT 28.6000 14.2000 28.9000 15.9000 ;
	    RECT 30.2500 15.2000 30.5500 21.8000 ;
	    RECT 31.7000 15.9000 32.1000 16.3000 ;
	    RECT 33.4500 16.2000 33.7500 25.8000 ;
	    RECT 35.8500 25.2000 36.1500 25.8000 ;
	    RECT 41.4500 25.2000 41.7500 25.8000 ;
	    RECT 35.8000 24.8000 36.2000 25.2000 ;
	    RECT 38.2000 25.1500 38.6000 25.2000 ;
	    RECT 39.0000 25.1500 39.4000 25.2000 ;
	    RECT 38.2000 24.8500 39.4000 25.1500 ;
	    RECT 38.2000 24.8000 38.6000 24.8500 ;
	    RECT 39.0000 24.8000 39.4000 24.8500 ;
	    RECT 41.4000 24.8000 41.8000 25.2000 ;
	    RECT 44.6000 25.1000 44.9000 26.8000 ;
	    RECT 45.4000 26.1500 45.8000 26.2000 ;
	    RECT 46.2000 26.1500 46.6000 26.2000 ;
	    RECT 45.4000 25.8500 46.6000 26.1500 ;
	    RECT 45.4000 25.8000 45.8000 25.8500 ;
	    RECT 46.2000 25.8000 46.6000 25.8500 ;
	    RECT 47.1000 26.1000 47.4000 26.8000 ;
	    RECT 47.1000 25.7000 47.5000 26.1000 ;
	    RECT 47.8000 25.1000 48.1000 27.5000 ;
	    RECT 52.6000 27.5000 53.0000 27.9000 ;
	    RECT 55.7000 27.8000 56.1000 27.9000 ;
	    RECT 53.3000 27.5000 56.1000 27.8000 ;
	    RECT 51.8000 26.8000 52.2000 27.2000 ;
	    RECT 52.6000 27.1000 52.9000 27.5000 ;
	    RECT 53.3000 27.4000 53.7000 27.5000 ;
	    RECT 55.0000 27.4000 55.4000 27.5000 ;
	    RECT 52.6000 26.8000 55.4000 27.1000 ;
	    RECT 51.8500 26.2000 52.1500 26.8000 ;
	    RECT 51.8000 25.8000 52.2000 26.2000 ;
	    RECT 44.6000 24.7000 45.0000 25.1000 ;
	    RECT 47.7000 24.7000 48.1000 25.1000 ;
	    RECT 52.6000 25.1000 52.9000 26.8000 ;
	    RECT 53.4000 26.1500 53.8000 26.2000 ;
	    RECT 54.2000 26.1500 54.6000 26.2000 ;
	    RECT 53.4000 25.8500 54.6000 26.1500 ;
	    RECT 53.4000 25.8000 53.8000 25.8500 ;
	    RECT 54.2000 25.8000 54.6000 25.8500 ;
	    RECT 55.1000 26.1000 55.4000 26.8000 ;
	    RECT 55.1000 25.7000 55.5000 26.1000 ;
	    RECT 55.8000 25.1000 56.1000 27.5000 ;
	    RECT 56.6000 26.8000 57.0000 27.2000 ;
	    RECT 52.6000 24.7000 53.0000 25.1000 ;
	    RECT 55.7000 24.7000 56.1000 25.1000 ;
	    RECT 39.8000 23.8000 40.2000 24.2000 ;
	    RECT 35.8000 21.8000 36.2000 22.2000 ;
	    RECT 30.2000 14.8000 30.6000 15.2000 ;
	    RECT 31.1000 14.9000 31.5000 15.3000 ;
	    RECT 31.1000 14.2000 31.4000 14.9000 ;
	    RECT 27.8000 13.8000 28.2000 14.2000 ;
	    RECT 28.6000 13.9000 31.4000 14.2000 ;
	    RECT 28.6000 13.5000 28.9000 13.9000 ;
	    RECT 29.3000 13.5000 29.7000 13.6000 ;
	    RECT 31.0000 13.5000 31.4000 13.6000 ;
	    RECT 31.8000 13.5000 32.1000 15.9000 ;
	    RECT 33.4000 15.8000 33.8000 16.2000 ;
	    RECT 33.4500 14.2000 33.7500 15.8000 ;
	    RECT 35.8500 14.2000 36.1500 21.8000 ;
	    RECT 39.0000 15.8000 39.4000 16.2000 ;
	    RECT 39.8500 16.1500 40.1500 23.8000 ;
	    RECT 56.6500 19.2000 56.9500 26.8000 ;
	    RECT 58.2000 25.8000 58.6000 26.2000 ;
	    RECT 61.4000 25.8000 61.8000 26.2000 ;
	    RECT 58.2500 25.2000 58.5500 25.8000 ;
	    RECT 58.2000 24.8000 58.6000 25.2000 ;
	    RECT 57.4000 21.8000 57.8000 22.2000 ;
	    RECT 53.4000 18.8000 53.8000 19.2000 ;
	    RECT 56.6000 18.8000 57.0000 19.2000 ;
	    RECT 42.2000 17.1500 42.6000 17.2000 ;
	    RECT 43.0000 17.1500 43.4000 17.2000 ;
	    RECT 42.2000 16.8500 43.4000 17.1500 ;
	    RECT 42.2000 16.8000 42.6000 16.8500 ;
	    RECT 43.0000 16.8000 43.4000 16.8500 ;
	    RECT 45.4000 16.8000 45.8000 17.2000 ;
	    RECT 45.4500 16.2000 45.7500 16.8000 ;
	    RECT 40.6000 16.1500 41.0000 16.2000 ;
	    RECT 39.8500 15.8500 41.0000 16.1500 ;
	    RECT 40.6000 15.8000 41.0000 15.8500 ;
	    RECT 42.2000 16.1500 42.6000 16.2000 ;
	    RECT 43.0000 16.1500 43.4000 16.2000 ;
	    RECT 42.2000 15.8500 43.4000 16.1500 ;
	    RECT 42.2000 15.8000 42.6000 15.8500 ;
	    RECT 43.0000 15.8000 43.4000 15.8500 ;
	    RECT 45.4000 15.8000 45.8000 16.2000 ;
	    RECT 39.0500 15.2000 39.3500 15.8000 ;
	    RECT 40.6500 15.2000 40.9500 15.8000 ;
	    RECT 39.0000 14.8000 39.4000 15.2000 ;
	    RECT 40.6000 14.8000 41.0000 15.2000 ;
	    RECT 43.0000 14.8000 43.4000 15.2000 ;
	    RECT 43.0500 14.2000 43.3500 14.8000 ;
	    RECT 53.4500 14.2000 53.7500 18.8000 ;
	    RECT 57.4500 17.2000 57.7500 21.8000 ;
	    RECT 57.4000 16.8000 57.8000 17.2000 ;
	    RECT 54.2000 15.8000 54.6000 16.2000 ;
	    RECT 57.4000 15.9000 57.8000 16.3000 ;
	    RECT 59.0000 16.1500 59.4000 16.2000 ;
	    RECT 59.8000 16.1500 60.2000 16.2000 ;
	    RECT 32.6000 13.8000 33.0000 14.2000 ;
	    RECT 33.4000 13.8000 33.8000 14.2000 ;
	    RECT 35.8000 13.8000 36.2000 14.2000 ;
	    RECT 39.0000 14.1500 39.4000 14.2000 ;
	    RECT 39.8000 14.1500 40.2000 14.2000 ;
	    RECT 39.0000 13.8500 40.2000 14.1500 ;
	    RECT 39.0000 13.8000 39.4000 13.8500 ;
	    RECT 39.8000 13.8000 40.2000 13.8500 ;
	    RECT 43.0000 13.8000 43.4000 14.2000 ;
	    RECT 44.6000 14.1500 45.0000 14.2000 ;
	    RECT 45.4000 14.1500 45.8000 14.2000 ;
	    RECT 44.6000 13.8500 45.8000 14.1500 ;
	    RECT 44.6000 13.8000 45.0000 13.8500 ;
	    RECT 45.4000 13.8000 45.8000 13.8500 ;
	    RECT 47.0000 14.1500 47.4000 14.2000 ;
	    RECT 47.8000 14.1500 48.2000 14.2000 ;
	    RECT 47.0000 13.8500 48.2000 14.1500 ;
	    RECT 47.0000 13.8000 47.4000 13.8500 ;
	    RECT 47.8000 13.8000 48.2000 13.8500 ;
	    RECT 52.6000 14.1500 53.0000 14.2000 ;
	    RECT 53.4000 14.1500 53.8000 14.2000 ;
	    RECT 52.6000 13.8500 53.8000 14.1500 ;
	    RECT 52.6000 13.8000 53.0000 13.8500 ;
	    RECT 53.4000 13.8000 53.8000 13.8500 ;
	    RECT 23.0000 12.8000 23.4000 13.2000 ;
	    RECT 23.8000 12.8000 24.2000 13.2000 ;
	    RECT 28.6000 13.1000 29.0000 13.5000 ;
	    RECT 29.3000 13.2000 32.1000 13.5000 ;
	    RECT 32.6500 13.2000 32.9500 13.8000 ;
	    RECT 35.8500 13.2000 36.1500 13.8000 ;
	    RECT 54.2500 13.2000 54.5500 15.8000 ;
	    RECT 57.4000 14.2000 57.7000 15.9000 ;
	    RECT 59.0000 15.8500 60.2000 16.1500 ;
	    RECT 60.5000 15.9000 60.9000 16.3000 ;
	    RECT 59.0000 15.8000 59.4000 15.8500 ;
	    RECT 59.8000 15.8000 60.2000 15.8500 ;
	    RECT 59.9000 14.9000 60.3000 15.3000 ;
	    RECT 59.9000 14.2000 60.2000 14.9000 ;
	    RECT 55.8000 13.8000 56.2000 14.2000 ;
	    RECT 56.6000 13.8000 57.0000 14.2000 ;
	    RECT 57.4000 13.9000 60.2000 14.2000 ;
	    RECT 31.7000 13.1000 32.1000 13.2000 ;
	    RECT 32.6000 12.8000 33.0000 13.2000 ;
	    RECT 35.8000 12.8000 36.2000 13.2000 ;
	    RECT 38.2000 13.1500 38.6000 13.2000 ;
	    RECT 39.0000 13.1500 39.4000 13.2000 ;
	    RECT 38.2000 12.8500 39.4000 13.1500 ;
	    RECT 38.2000 12.8000 38.6000 12.8500 ;
	    RECT 39.0000 12.8000 39.4000 12.8500 ;
	    RECT 43.0000 12.8000 43.4000 13.2000 ;
	    RECT 50.2000 12.8000 50.6000 13.2000 ;
	    RECT 54.2000 12.8000 54.6000 13.2000 ;
	    RECT 23.8500 12.2000 24.1500 12.8000 ;
	    RECT 23.8000 11.8000 24.2000 12.2000 ;
	    RECT 26.2000 11.8000 26.6000 12.2000 ;
	    RECT 30.2000 11.8000 30.6000 12.2000 ;
	    RECT 33.4000 11.8000 33.8000 12.2000 ;
	    RECT 36.6000 11.8000 37.0000 12.2000 ;
	    RECT 19.8000 8.8000 20.2000 9.2000 ;
	    RECT 21.4000 8.8000 21.8000 9.2000 ;
	    RECT 22.2000 9.1500 22.6000 9.2000 ;
	    RECT 23.0000 9.1500 23.4000 9.2000 ;
	    RECT 22.2000 8.8500 23.4000 9.1500 ;
	    RECT 22.2000 8.8000 22.6000 8.8500 ;
	    RECT 23.0000 8.8000 23.4000 8.8500 ;
	    RECT 26.2500 8.2000 26.5500 11.8000 ;
	    RECT 29.4000 8.8000 29.8000 9.2000 ;
	    RECT 29.4500 8.2000 29.7500 8.8000 ;
	    RECT 22.2000 7.8000 22.6000 8.2000 ;
	    RECT 26.2000 7.8000 26.6000 8.2000 ;
	    RECT 29.4000 7.8000 29.8000 8.2000 ;
	    RECT 22.2500 7.2000 22.5500 7.8000 ;
	    RECT 22.2000 7.1500 22.6000 7.2000 ;
	    RECT 23.0000 7.1500 23.4000 7.2000 ;
	    RECT 30.2500 7.1500 30.5500 11.8000 ;
	    RECT 22.2000 6.8500 23.4000 7.1500 ;
	    RECT 22.2000 6.8000 22.6000 6.8500 ;
	    RECT 23.0000 6.8000 23.4000 6.8500 ;
	    RECT 29.4500 6.8500 30.5500 7.1500 ;
	    RECT 29.4500 6.2000 29.7500 6.8500 ;
	    RECT 15.8000 6.1500 16.2000 6.2000 ;
	    RECT 15.0500 5.8500 16.2000 6.1500 ;
	    RECT 15.0500 5.2000 15.3500 5.8500 ;
	    RECT 15.8000 5.8000 16.2000 5.8500 ;
	    RECT 29.4000 5.8000 29.8000 6.2000 ;
	    RECT 33.4500 5.2000 33.7500 11.8000 ;
	    RECT 35.8000 7.8000 36.2000 8.2000 ;
	    RECT 35.8500 7.2000 36.1500 7.8000 ;
	    RECT 35.8000 6.8000 36.2000 7.2000 ;
	    RECT 36.6500 5.2000 36.9500 11.8000 ;
	    RECT 43.0500 9.2000 43.3500 12.8000 ;
	    RECT 45.4000 12.1500 45.8000 12.2000 ;
	    RECT 46.2000 12.1500 46.6000 12.2000 ;
	    RECT 45.4000 11.8500 46.6000 12.1500 ;
	    RECT 45.4000 11.8000 45.8000 11.8500 ;
	    RECT 46.2000 11.8000 46.6000 11.8500 ;
	    RECT 50.2500 9.2000 50.5500 12.8000 ;
	    RECT 51.0000 11.8000 51.4000 12.2000 ;
	    RECT 51.0500 9.2000 51.3500 11.8000 ;
	    RECT 55.8500 9.2000 56.1500 13.8000 ;
	    RECT 56.6500 12.2000 56.9500 13.8000 ;
	    RECT 57.4000 13.5000 57.7000 13.9000 ;
	    RECT 58.1000 13.5000 58.5000 13.6000 ;
	    RECT 59.8000 13.5000 60.2000 13.6000 ;
	    RECT 60.6000 13.5000 60.9000 15.9000 ;
	    RECT 61.4500 15.2000 61.7500 25.8000 ;
	    RECT 62.2000 15.8000 62.6000 16.2000 ;
	    RECT 62.2500 15.2000 62.5500 15.8000 ;
	    RECT 61.4000 14.8000 61.8000 15.2000 ;
	    RECT 62.2000 14.8000 62.6000 15.2000 ;
	    RECT 61.4000 13.8000 61.8000 14.2000 ;
	    RECT 57.4000 13.1000 57.8000 13.5000 ;
	    RECT 58.1000 13.2000 60.9000 13.5000 ;
	    RECT 61.4500 13.2000 61.7500 13.8000 ;
	    RECT 60.5000 13.1000 60.9000 13.2000 ;
	    RECT 61.4000 12.8000 61.8000 13.2000 ;
	    RECT 56.6000 11.8000 57.0000 12.2000 ;
	    RECT 39.8000 9.1500 40.2000 9.2000 ;
	    RECT 40.6000 9.1500 41.0000 9.2000 ;
	    RECT 39.8000 8.8500 41.0000 9.1500 ;
	    RECT 39.8000 8.8000 40.2000 8.8500 ;
	    RECT 40.6000 8.8000 41.0000 8.8500 ;
	    RECT 43.0000 8.8000 43.4000 9.2000 ;
	    RECT 50.2000 8.8000 50.6000 9.2000 ;
	    RECT 51.0000 8.8000 51.4000 9.2000 ;
	    RECT 55.8000 8.8000 56.2000 9.2000 ;
	    RECT 59.8000 9.1500 60.2000 9.2000 ;
	    RECT 60.6000 9.1500 61.0000 9.2000 ;
	    RECT 59.8000 8.8500 61.0000 9.1500 ;
	    RECT 59.8000 8.8000 60.2000 8.8500 ;
	    RECT 60.6000 8.8000 61.0000 8.8500 ;
	    RECT 48.6000 7.5000 49.0000 7.9000 ;
	    RECT 51.7000 7.8000 52.1000 7.9000 ;
	    RECT 49.3000 7.5000 52.1000 7.8000 ;
	    RECT 39.0000 6.8000 39.4000 7.2000 ;
	    RECT 40.6000 7.1500 41.0000 7.2000 ;
	    RECT 41.4000 7.1500 41.8000 7.2000 ;
	    RECT 40.6000 6.8500 41.8000 7.1500 ;
	    RECT 40.6000 6.8000 41.0000 6.8500 ;
	    RECT 41.4000 6.8000 41.8000 6.8500 ;
	    RECT 43.0000 6.8000 43.4000 7.2000 ;
	    RECT 48.6000 7.1000 48.9000 7.5000 ;
	    RECT 49.3000 7.4000 49.7000 7.5000 ;
	    RECT 51.0000 7.4000 51.4000 7.5000 ;
	    RECT 48.6000 6.8000 51.4000 7.1000 ;
	    RECT 39.0500 6.2000 39.3500 6.8000 ;
	    RECT 43.0500 6.2000 43.3500 6.8000 ;
	    RECT 39.0000 5.8000 39.4000 6.2000 ;
	    RECT 40.6000 6.1500 41.0000 6.2000 ;
	    RECT 41.4000 6.1500 41.8000 6.2000 ;
	    RECT 40.6000 5.8500 41.8000 6.1500 ;
	    RECT 40.6000 5.8000 41.0000 5.8500 ;
	    RECT 41.4000 5.8000 41.8000 5.8500 ;
	    RECT 43.0000 5.8000 43.4000 6.2000 ;
	    RECT 3.8000 4.7000 4.2000 5.1000 ;
	    RECT 6.9000 4.7000 7.3000 5.1000 ;
	    RECT 10.2000 5.1500 10.6000 5.2000 ;
	    RECT 11.0000 5.1500 11.4000 5.2000 ;
	    RECT 10.2000 4.8500 11.4000 5.1500 ;
	    RECT 10.2000 4.8000 10.6000 4.8500 ;
	    RECT 11.0000 4.8000 11.4000 4.8500 ;
	    RECT 15.0000 4.8000 15.4000 5.2000 ;
	    RECT 33.4000 4.8000 33.8000 5.2000 ;
	    RECT 36.6000 4.8000 37.0000 5.2000 ;
	    RECT 48.6000 5.1000 48.9000 6.8000 ;
	    RECT 51.1000 6.1000 51.4000 6.8000 ;
	    RECT 51.1000 5.7000 51.5000 6.1000 ;
	    RECT 51.8000 5.1000 52.1000 7.5000 ;
	    RECT 58.3000 7.8000 58.7000 7.9000 ;
	    RECT 58.3000 7.5000 61.1000 7.8000 ;
	    RECT 61.4000 7.5000 61.8000 7.9000 ;
	    RECT 55.8000 6.1500 56.2000 6.2000 ;
	    RECT 56.6000 6.1500 57.0000 6.2000 ;
	    RECT 55.8000 5.8500 57.0000 6.1500 ;
	    RECT 55.8000 5.8000 56.2000 5.8500 ;
	    RECT 56.6000 5.8000 57.0000 5.8500 ;
	    RECT 48.6000 4.7000 49.0000 5.1000 ;
	    RECT 51.7000 4.7000 52.1000 5.1000 ;
	    RECT 58.3000 5.1000 58.6000 7.5000 ;
	    RECT 59.0000 7.4000 59.4000 7.5000 ;
	    RECT 60.7000 7.4000 61.1000 7.5000 ;
	    RECT 61.5000 7.1000 61.8000 7.5000 ;
	    RECT 59.0000 6.8000 61.8000 7.1000 ;
	    RECT 59.0000 6.1000 59.3000 6.8000 ;
	    RECT 58.9000 5.7000 59.3000 6.1000 ;
	    RECT 61.5000 5.1000 61.8000 6.8000 ;
	    RECT 58.3000 4.7000 58.7000 5.1000 ;
	    RECT 61.4000 4.7000 61.8000 5.1000 ;
         LAYER metal3 ;
	    RECT 7.8000 29.1500 8.2000 29.2000 ;
	    RECT 11.0000 29.1500 11.4000 29.2000 ;
	    RECT 7.8000 28.8500 11.4000 29.1500 ;
	    RECT 7.8000 28.8000 8.2000 28.8500 ;
	    RECT 11.0000 28.8000 11.4000 28.8500 ;
	    RECT 38.2000 28.1500 38.6000 28.2000 ;
	    RECT 39.8000 28.1500 40.2000 28.2000 ;
	    RECT 38.2000 27.8500 40.2000 28.1500 ;
	    RECT 38.2000 27.8000 38.6000 27.8500 ;
	    RECT 39.8000 27.8000 40.2000 27.8500 ;
	    RECT 29.4000 27.1500 29.8000 27.2000 ;
	    RECT 34.2000 27.1500 34.6000 27.2000 ;
	    RECT 29.4000 26.8500 34.6000 27.1500 ;
	    RECT 29.4000 26.8000 29.8000 26.8500 ;
	    RECT 34.2000 26.8000 34.6000 26.8500 ;
	    RECT 1.4000 26.1500 1.8000 26.2000 ;
	    RECT 46.2000 26.1500 46.6000 26.2000 ;
	    RECT 51.8000 26.1500 52.2000 26.2000 ;
	    RECT 1.4000 25.8500 5.7500 26.1500 ;
	    RECT 1.4000 25.8000 1.8000 25.8500 ;
	    RECT 5.4500 25.2000 5.7500 25.8500 ;
	    RECT 46.2000 25.8500 52.2000 26.1500 ;
	    RECT 46.2000 25.8000 46.6000 25.8500 ;
	    RECT 51.8000 25.8000 52.2000 25.8500 ;
	    RECT 53.4000 26.1500 53.8000 26.2000 ;
	    RECT 58.2000 26.1500 58.6000 26.2000 ;
	    RECT 53.4000 25.8500 58.6000 26.1500 ;
	    RECT 53.4000 25.8000 53.8000 25.8500 ;
	    RECT 58.2000 25.8000 58.6000 25.8500 ;
	    RECT 3.0000 25.1500 3.4000 25.2000 ;
	    RECT 3.8000 25.1500 4.2000 25.2000 ;
	    RECT 3.0000 24.8500 4.2000 25.1500 ;
	    RECT 3.0000 24.8000 3.4000 24.8500 ;
	    RECT 3.8000 24.8000 4.2000 24.8500 ;
	    RECT 5.4000 24.8000 5.8000 25.2000 ;
	    RECT 35.8000 25.1500 36.2000 25.2000 ;
	    RECT 39.0000 25.1500 39.4000 25.2000 ;
	    RECT 41.4000 25.1500 41.8000 25.2000 ;
	    RECT 35.8000 24.8500 41.8000 25.1500 ;
	    RECT 35.8000 24.8000 36.2000 24.8500 ;
	    RECT 39.0000 24.8000 39.4000 24.8500 ;
	    RECT 41.4000 24.8000 41.8000 24.8500 ;
	    RECT 19.0000 22.1500 19.4000 22.2000 ;
	    RECT 20.6000 22.1500 21.0000 22.2000 ;
	    RECT 19.0000 21.8500 21.0000 22.1500 ;
	    RECT 19.0000 21.8000 19.4000 21.8500 ;
	    RECT 20.6000 21.8000 21.0000 21.8500 ;
	    RECT 24.6000 22.1500 25.0000 22.2000 ;
	    RECT 27.8000 22.1500 28.2000 22.2000 ;
	    RECT 24.6000 21.8500 28.2000 22.1500 ;
	    RECT 24.6000 21.8000 25.0000 21.8500 ;
	    RECT 27.8000 21.8000 28.2000 21.8500 ;
	    RECT 53.4000 19.1500 53.8000 19.2000 ;
	    RECT 56.6000 19.1500 57.0000 19.2000 ;
	    RECT 53.4000 18.8500 57.0000 19.1500 ;
	    RECT 53.4000 18.8000 53.8000 18.8500 ;
	    RECT 56.6000 18.8000 57.0000 18.8500 ;
	    RECT 22.2000 16.8000 22.6000 17.2000 ;
	    RECT 43.0000 17.1500 43.4000 17.2000 ;
	    RECT 45.4000 17.1500 45.8000 17.2000 ;
	    RECT 42.2500 16.8500 45.8000 17.1500 ;
	    RECT 43.0000 16.8000 43.4000 16.8500 ;
	    RECT 45.4000 16.8000 45.8000 16.8500 ;
	    RECT 56.6000 17.1500 57.0000 17.2000 ;
	    RECT 57.4000 17.1500 57.8000 17.2000 ;
	    RECT 56.6000 16.8500 57.8000 17.1500 ;
	    RECT 56.6000 16.8000 57.0000 16.8500 ;
	    RECT 57.4000 16.8000 57.8000 16.8500 ;
	    RECT 22.2500 16.1500 22.5500 16.8000 ;
	    RECT 26.2000 16.1500 26.6000 16.2000 ;
	    RECT 22.2500 15.8500 26.6000 16.1500 ;
	    RECT 26.2000 15.8000 26.6000 15.8500 ;
	    RECT 40.6000 16.1500 41.0000 16.2000 ;
	    RECT 42.2000 16.1500 42.6000 16.2000 ;
	    RECT 40.6000 15.8500 42.6000 16.1500 ;
	    RECT 40.6000 15.8000 41.0000 15.8500 ;
	    RECT 42.2000 15.8000 42.6000 15.8500 ;
	    RECT 59.8000 16.1500 60.2000 16.2000 ;
	    RECT 62.2000 16.1500 62.6000 16.2000 ;
	    RECT 59.8000 15.8500 62.6000 16.1500 ;
	    RECT 59.8000 15.8000 60.2000 15.8500 ;
	    RECT 62.2000 15.8000 62.6000 15.8500 ;
	    RECT 7.8000 15.1500 8.2000 15.2000 ;
	    RECT 8.6000 15.1500 9.0000 15.2000 ;
	    RECT 13.4000 15.1500 13.8000 15.2000 ;
	    RECT 7.8000 14.8500 13.8000 15.1500 ;
	    RECT 7.8000 14.8000 8.2000 14.8500 ;
	    RECT 8.6000 14.8000 9.0000 14.8500 ;
	    RECT 13.4000 14.8000 13.8000 14.8500 ;
	    RECT 14.2000 15.1500 14.6000 15.2000 ;
	    RECT 18.2000 15.1500 18.6000 15.2000 ;
	    RECT 14.2000 14.8500 18.6000 15.1500 ;
	    RECT 14.2000 14.8000 14.6000 14.8500 ;
	    RECT 18.2000 14.8000 18.6000 14.8500 ;
	    RECT 29.4000 15.1500 29.8000 15.2000 ;
	    RECT 30.2000 15.1500 30.6000 15.2000 ;
	    RECT 29.4000 14.8500 30.6000 15.1500 ;
	    RECT 29.4000 14.8000 29.8000 14.8500 ;
	    RECT 30.2000 14.8000 30.6000 14.8500 ;
	    RECT 39.0000 15.1500 39.4000 15.2000 ;
	    RECT 43.0000 15.1500 43.4000 15.2000 ;
	    RECT 39.0000 14.8500 43.4000 15.1500 ;
	    RECT 39.0000 14.8000 39.4000 14.8500 ;
	    RECT 43.0000 14.8000 43.4000 14.8500 ;
	    RECT 59.8000 15.1500 60.2000 15.2000 ;
	    RECT 61.4000 15.1500 61.8000 15.2000 ;
	    RECT 59.8000 14.8500 61.8000 15.1500 ;
	    RECT 59.8000 14.8000 60.2000 14.8500 ;
	    RECT 61.4000 14.8000 61.8000 14.8500 ;
	    RECT 16.6000 14.1500 17.0000 14.2000 ;
	    RECT 20.6000 14.1500 21.0000 14.2000 ;
	    RECT 16.6000 13.8500 21.0000 14.1500 ;
	    RECT 16.6000 13.8000 17.0000 13.8500 ;
	    RECT 20.6000 13.8000 21.0000 13.8500 ;
	    RECT 33.4000 14.1500 33.8000 14.2000 ;
	    RECT 39.0000 14.1500 39.4000 14.2000 ;
	    RECT 33.4000 13.8500 39.4000 14.1500 ;
	    RECT 33.4000 13.8000 33.8000 13.8500 ;
	    RECT 39.0000 13.8000 39.4000 13.8500 ;
	    RECT 45.4000 14.1500 45.8000 14.2000 ;
	    RECT 47.8000 14.1500 48.2000 14.2000 ;
	    RECT 52.6000 14.1500 53.0000 14.2000 ;
	    RECT 45.4000 13.8500 53.0000 14.1500 ;
	    RECT 45.4000 13.8000 45.8000 13.8500 ;
	    RECT 47.8000 13.8000 48.2000 13.8500 ;
	    RECT 52.6000 13.8000 53.0000 13.8500 ;
	    RECT 55.8000 14.1500 56.2000 14.2000 ;
	    RECT 55.8000 13.8500 61.7500 14.1500 ;
	    RECT 55.8000 13.8000 56.2000 13.8500 ;
	    RECT 61.4500 13.2000 61.7500 13.8500 ;
	    RECT 9.4000 13.1500 9.8000 13.2000 ;
	    RECT 10.2000 13.1500 10.6000 13.2000 ;
	    RECT 9.4000 12.8500 10.6000 13.1500 ;
	    RECT 9.4000 12.8000 9.8000 12.8500 ;
	    RECT 10.2000 12.8000 10.6000 12.8500 ;
	    RECT 13.4000 13.1500 13.8000 13.2000 ;
	    RECT 23.0000 13.1500 23.4000 13.2000 ;
	    RECT 13.4000 12.8500 23.4000 13.1500 ;
	    RECT 13.4000 12.8000 13.8000 12.8500 ;
	    RECT 23.0000 12.8000 23.4000 12.8500 ;
	    RECT 32.6000 13.1500 33.0000 13.2000 ;
	    RECT 39.0000 13.1500 39.4000 13.2000 ;
	    RECT 32.6000 12.8500 39.4000 13.1500 ;
	    RECT 32.6000 12.8000 33.0000 12.8500 ;
	    RECT 39.0000 12.8000 39.4000 12.8500 ;
	    RECT 43.0000 13.1500 43.4000 13.2000 ;
	    RECT 54.2000 13.1500 54.6000 13.2000 ;
	    RECT 43.0000 12.8500 54.6000 13.1500 ;
	    RECT 43.0000 12.8000 43.4000 12.8500 ;
	    RECT 54.2000 12.8000 54.6000 12.8500 ;
	    RECT 61.4000 12.8000 61.8000 13.2000 ;
	    RECT 11.0000 12.1500 11.4000 12.2000 ;
	    RECT 23.8000 12.1500 24.2000 12.2000 ;
	    RECT 10.2500 11.8500 24.2000 12.1500 ;
	    RECT 11.0000 11.8000 11.4000 11.8500 ;
	    RECT 23.8000 11.8000 24.2000 11.8500 ;
	    RECT 36.6000 12.1500 37.0000 12.2000 ;
	    RECT 46.2000 12.1500 46.6000 12.2000 ;
	    RECT 36.6000 11.8500 46.6000 12.1500 ;
	    RECT 36.6000 11.8000 37.0000 11.8500 ;
	    RECT 46.2000 11.8000 46.6000 11.8500 ;
	    RECT 51.0000 12.1500 51.4000 12.2000 ;
	    RECT 56.6000 12.1500 57.0000 12.2000 ;
	    RECT 51.0000 11.8500 57.0000 12.1500 ;
	    RECT 51.0000 11.8000 51.4000 11.8500 ;
	    RECT 56.6000 11.8000 57.0000 11.8500 ;
	    RECT 14.2000 9.1500 14.6000 9.2000 ;
	    RECT 19.8000 9.1500 20.2000 9.2000 ;
	    RECT 14.2000 8.8500 20.2000 9.1500 ;
	    RECT 14.2000 8.8000 14.6000 8.8500 ;
	    RECT 19.8000 8.8000 20.2000 8.8500 ;
	    RECT 21.4000 9.1500 21.8000 9.2000 ;
	    RECT 22.2000 9.1500 22.6000 9.2000 ;
	    RECT 21.4000 8.8500 22.6000 9.1500 ;
	    RECT 21.4000 8.8000 21.8000 8.8500 ;
	    RECT 22.2000 8.8000 22.6000 8.8500 ;
	    RECT 29.4000 8.8000 29.8000 9.2000 ;
	    RECT 40.6000 9.1500 41.0000 9.2000 ;
	    RECT 50.2000 9.1500 50.6000 9.2000 ;
	    RECT 39.8500 8.8500 50.6000 9.1500 ;
	    RECT 40.6000 8.8000 41.0000 8.8500 ;
	    RECT 50.2000 8.8000 50.6000 8.8500 ;
	    RECT 59.8000 9.1500 60.2000 9.2000 ;
	    RECT 60.6000 9.1500 61.0000 9.2000 ;
	    RECT 59.8000 8.8500 61.0000 9.1500 ;
	    RECT 59.8000 8.8000 60.2000 8.8500 ;
	    RECT 60.6000 8.8000 61.0000 8.8500 ;
	    RECT 29.4500 8.2000 29.7500 8.8000 ;
	    RECT 3.0000 8.1500 3.4000 8.2000 ;
	    RECT 8.6000 8.1500 9.0000 8.2000 ;
	    RECT 22.2000 8.1500 22.6000 8.2000 ;
	    RECT 3.0000 7.8500 22.6000 8.1500 ;
	    RECT 3.0000 7.8000 3.4000 7.8500 ;
	    RECT 8.6000 7.8000 9.0000 7.8500 ;
	    RECT 22.2000 7.8000 22.6000 7.8500 ;
	    RECT 29.4000 7.8000 29.8000 8.2000 ;
	    RECT 35.8000 7.8000 36.2000 8.2000 ;
	    RECT 10.2000 7.1500 10.6000 7.2000 ;
	    RECT 7.8500 6.8500 10.6000 7.1500 ;
	    RECT 7.8500 6.2000 8.1500 6.8500 ;
	    RECT 10.2000 6.8000 10.6000 6.8500 ;
	    RECT 23.0000 7.1500 23.4000 7.2000 ;
	    RECT 35.8500 7.1500 36.1500 7.8000 ;
	    RECT 23.0000 6.8500 36.1500 7.1500 ;
	    RECT 39.0000 7.1500 39.4000 7.2000 ;
	    RECT 40.6000 7.1500 41.0000 7.2000 ;
	    RECT 39.0000 6.8500 41.0000 7.1500 ;
	    RECT 23.0000 6.8000 23.4000 6.8500 ;
	    RECT 39.0000 6.8000 39.4000 6.8500 ;
	    RECT 40.6000 6.8000 41.0000 6.8500 ;
	    RECT 7.8000 5.8000 8.2000 6.2000 ;
	    RECT 41.4000 6.1500 41.8000 6.2000 ;
	    RECT 43.0000 6.1500 43.4000 6.2000 ;
	    RECT 41.4000 5.8500 43.4000 6.1500 ;
	    RECT 41.4000 5.8000 41.8000 5.8500 ;
	    RECT 43.0000 5.8000 43.4000 5.8500 ;
	    RECT 55.8000 6.1500 56.2000 6.2000 ;
	    RECT 56.6000 6.1500 57.0000 6.2000 ;
	    RECT 55.8000 5.8500 57.0000 6.1500 ;
	    RECT 55.8000 5.8000 56.2000 5.8500 ;
	    RECT 56.6000 5.8000 57.0000 5.8500 ;
	    RECT 11.0000 5.1500 11.4000 5.2000 ;
	    RECT 15.0000 5.1500 15.4000 5.2000 ;
	    RECT 11.0000 4.8500 15.4000 5.1500 ;
	    RECT 11.0000 4.8000 11.4000 4.8500 ;
	    RECT 15.0000 4.8000 15.4000 4.8500 ;
         LAYER metal4 ;
	    RECT 3.8000 25.1500 4.2000 25.2000 ;
	    RECT 3.0500 24.8500 4.2000 25.1500 ;
	    RECT 3.0500 8.2000 3.3500 24.8500 ;
	    RECT 3.8000 24.8000 4.2000 24.8500 ;
	    RECT 56.6000 16.8000 57.0000 17.2000 ;
	    RECT 29.4000 14.8000 29.8000 15.2000 ;
	    RECT 29.4500 8.2000 29.7500 14.8000 ;
	    RECT 3.0000 7.8000 3.4000 8.2000 ;
	    RECT 29.4000 7.8000 29.8000 8.2000 ;
	    RECT 56.6500 6.2000 56.9500 16.8000 ;
	    RECT 59.8000 14.8000 60.2000 15.2000 ;
	    RECT 59.8500 9.2000 60.1500 14.8000 ;
	    RECT 59.8000 8.8000 60.2000 9.2000 ;
	    RECT 56.6000 5.8000 57.0000 6.2000 ;
   END
END adder
