magic
tech scmos
magscale 1 2
timestamp 1591289005
<< metal1 >>
rect 938 614 950 616
rect 928 606 930 614
rect 938 606 940 614
rect 948 606 950 614
rect 958 606 960 614
rect 938 604 950 606
rect 212 576 216 584
rect 573 557 595 563
rect 285 543 291 556
rect 269 537 291 543
rect 573 537 595 543
rect 589 524 595 537
rect 861 543 867 563
rect 804 537 819 543
rect 861 537 876 543
rect 621 517 659 523
rect 676 517 691 523
rect 916 517 931 523
rect 1165 517 1187 523
rect 653 497 675 503
rect 829 503 835 516
rect 1165 504 1171 517
rect 829 497 851 503
rect 292 477 307 483
rect 781 477 796 483
rect 1261 477 1292 483
rect 333 437 364 443
rect 500 436 508 444
rect 612 436 614 444
rect 346 414 358 416
rect 336 406 338 414
rect 346 406 348 414
rect 356 406 358 414
rect 366 406 368 414
rect 346 404 358 406
rect 157 303 163 316
rect 141 297 163 303
rect 1069 303 1075 323
rect 861 297 883 303
rect 1069 297 1107 303
rect 861 284 867 297
rect 221 277 243 283
rect 189 263 195 276
rect 221 264 227 277
rect 397 277 435 283
rect 493 277 515 283
rect 701 277 716 283
rect 733 277 755 283
rect 1021 277 1043 283
rect 1053 277 1068 283
rect 1277 277 1292 283
rect 173 257 195 263
rect 298 236 300 244
rect 532 236 534 244
rect 938 214 950 216
rect 928 206 930 214
rect 938 206 940 214
rect 948 206 950 214
rect 958 206 960 214
rect 938 204 950 206
rect 1016 176 1020 184
rect 644 157 675 163
rect 228 137 243 143
rect 253 137 275 143
rect 292 137 307 143
rect 493 137 515 143
rect 605 137 627 143
rect 685 137 707 143
rect 781 143 787 163
rect 893 157 947 163
rect 749 137 787 143
rect 781 124 787 137
rect 941 143 947 157
rect 941 137 963 143
rect 45 117 115 123
rect 189 117 227 123
rect 221 97 227 117
rect 573 117 588 123
rect 861 123 867 136
rect 957 123 963 137
rect 1101 143 1107 163
rect 1069 137 1107 143
rect 1245 137 1260 143
rect 861 117 883 123
rect 957 117 988 123
rect 349 97 419 103
rect 429 97 467 103
rect 653 97 668 103
rect 861 97 883 103
rect 346 14 358 16
rect 336 6 338 14
rect 346 6 348 14
rect 356 6 358 14
rect 366 6 368 14
rect 346 4 358 6
<< m2contact >>
rect 920 606 928 614
rect 930 606 938 614
rect 940 606 948 614
rect 950 606 958 614
rect 960 606 968 614
rect 204 576 212 584
rect 396 576 404 584
rect 1212 576 1220 584
rect 284 556 292 564
rect 316 556 324 564
rect 556 556 564 564
rect 636 556 644 564
rect 748 556 756 564
rect 828 556 836 564
rect 60 536 68 544
rect 156 536 164 544
rect 172 536 180 544
rect 444 536 452 544
rect 540 536 548 544
rect 700 536 708 544
rect 796 536 804 544
rect 1164 556 1172 564
rect 876 536 884 544
rect 972 536 980 544
rect 1036 536 1044 544
rect 1132 536 1140 544
rect 44 516 52 524
rect 108 516 116 524
rect 428 516 436 524
rect 588 516 596 524
rect 668 516 676 524
rect 716 516 724 524
rect 828 516 836 524
rect 908 516 916 524
rect 1084 516 1092 524
rect 764 496 772 504
rect 1228 516 1236 524
rect 1164 496 1172 504
rect 12 476 20 484
rect 284 476 292 484
rect 796 476 804 484
rect 1292 476 1300 484
rect 364 436 372 444
rect 508 436 516 444
rect 604 436 612 444
rect 716 436 724 444
rect 1148 436 1156 444
rect 328 406 336 414
rect 338 406 346 414
rect 348 406 356 414
rect 358 406 366 414
rect 368 406 376 414
rect 844 336 852 344
rect 156 316 164 324
rect 268 316 276 324
rect 284 316 292 324
rect 444 316 452 324
rect 460 316 468 324
rect 540 316 548 324
rect 668 316 676 324
rect 780 316 788 324
rect 860 316 868 324
rect 908 316 916 324
rect 188 296 196 304
rect 380 296 388 304
rect 812 296 820 304
rect 1084 316 1092 324
rect 1180 316 1188 324
rect 1244 296 1252 304
rect 12 276 20 284
rect 108 276 116 284
rect 188 276 196 284
rect 124 256 132 264
rect 156 256 164 264
rect 316 276 324 284
rect 556 276 564 284
rect 652 276 660 284
rect 716 276 724 284
rect 796 276 804 284
rect 860 276 868 284
rect 892 276 900 284
rect 940 276 948 284
rect 1068 276 1076 284
rect 1116 276 1124 284
rect 1132 276 1140 284
rect 1228 276 1236 284
rect 1292 276 1300 284
rect 220 256 228 264
rect 412 256 420 264
rect 476 256 484 264
rect 716 256 724 264
rect 764 256 772 264
rect 1004 256 1012 264
rect 60 236 68 244
rect 204 236 212 244
rect 268 236 276 244
rect 300 236 308 244
rect 396 236 404 244
rect 524 236 532 244
rect 604 236 612 244
rect 668 236 676 244
rect 908 236 916 244
rect 920 206 928 214
rect 930 206 938 214
rect 940 206 948 214
rect 950 206 958 214
rect 960 206 968 214
rect 460 176 468 184
rect 796 176 804 184
rect 860 176 868 184
rect 1020 176 1028 184
rect 1116 176 1124 184
rect 1196 176 1204 184
rect 284 156 292 164
rect 524 156 532 164
rect 588 156 596 164
rect 764 156 772 164
rect 60 136 68 144
rect 156 136 164 144
rect 172 136 180 144
rect 220 136 228 144
rect 284 136 292 144
rect 444 136 452 144
rect 716 136 724 144
rect 828 136 836 144
rect 860 136 868 144
rect 1084 156 1092 164
rect 204 96 212 104
rect 316 116 324 124
rect 588 116 596 124
rect 780 116 788 124
rect 812 116 820 124
rect 1052 136 1060 144
rect 1148 136 1156 144
rect 1260 136 1268 144
rect 988 116 996 124
rect 1132 116 1140 124
rect 668 96 676 104
rect 732 96 740 104
rect 12 76 20 84
rect 540 36 548 44
rect 328 6 336 14
rect 338 6 346 14
rect 348 6 356 14
rect 358 6 366 14
rect 368 6 376 14
<< metal2 >>
rect 157 544 163 576
rect 173 544 179 616
rect 212 577 220 583
rect 285 564 291 683
rect 397 624 403 683
rect 317 564 323 616
rect 429 604 435 683
rect 397 584 403 596
rect 557 564 563 683
rect 637 564 643 683
rect 829 564 835 683
rect 756 557 764 563
rect 445 544 451 556
rect 541 544 547 556
rect 557 544 563 556
rect 797 544 803 556
rect 829 544 835 556
rect 877 544 883 683
rect 1197 677 1219 683
rect 938 614 950 616
rect 928 606 930 614
rect 938 606 940 614
rect 948 606 950 614
rect 958 606 960 614
rect 938 604 950 606
rect 1213 584 1219 677
rect 973 544 979 556
rect 692 537 700 543
rect 1165 543 1171 556
rect 1165 537 1187 543
rect 36 517 44 523
rect 61 504 67 536
rect 589 524 595 536
rect 1037 524 1043 536
rect 916 517 924 523
rect 1076 517 1084 523
rect 109 504 115 516
rect 13 484 19 496
rect 285 324 291 476
rect 372 437 380 443
rect 346 414 358 416
rect 336 406 338 414
rect 346 406 348 414
rect 356 406 358 414
rect 366 406 368 414
rect 346 404 358 406
rect 109 284 115 316
rect 157 304 163 316
rect 269 304 275 316
rect 285 304 291 316
rect 180 297 188 303
rect 372 297 380 303
rect 413 284 419 436
rect 116 277 124 283
rect 324 277 332 283
rect 13 264 19 276
rect 157 264 163 276
rect 189 264 195 276
rect 413 264 419 276
rect 132 257 140 263
rect 212 257 220 263
rect 269 244 275 256
rect 212 237 220 243
rect 61 144 67 236
rect 173 144 179 156
rect 212 137 220 143
rect 269 143 275 236
rect 285 164 291 176
rect 269 137 284 143
rect 157 124 163 136
rect 301 123 307 236
rect 397 184 403 236
rect 429 184 435 516
rect 500 437 508 443
rect 445 324 451 336
rect 532 317 540 323
rect 461 264 467 316
rect 557 284 563 436
rect 605 304 611 436
rect 669 324 675 516
rect 717 504 723 516
rect 829 504 835 516
rect 772 497 780 503
rect 669 284 675 316
rect 717 284 723 436
rect 797 323 803 476
rect 1133 384 1139 536
rect 1165 504 1171 516
rect 852 337 860 343
rect 909 324 915 336
rect 797 317 812 323
rect 852 317 860 323
rect 781 304 787 316
rect 813 304 819 316
rect 861 284 867 296
rect 1069 284 1075 376
rect 1149 344 1155 436
rect 1181 364 1187 537
rect 1188 317 1196 323
rect 788 277 796 283
rect 900 277 908 283
rect 948 277 956 283
rect 1060 277 1068 283
rect 653 264 659 276
rect 717 264 723 276
rect 1085 264 1091 316
rect 1229 304 1235 516
rect 1293 484 1299 496
rect 1245 304 1251 316
rect 772 257 780 263
rect 477 244 483 256
rect 452 177 460 183
rect 525 164 531 236
rect 589 164 595 176
rect 445 144 451 156
rect 452 137 460 143
rect 605 143 611 236
rect 589 137 611 143
rect 589 124 595 137
rect 301 117 316 123
rect 301 104 307 117
rect 669 104 675 236
rect 717 144 723 156
rect 733 104 739 236
rect 861 184 867 256
rect 916 237 924 243
rect 938 214 950 216
rect 928 206 930 214
rect 938 206 940 214
rect 948 206 950 214
rect 958 206 960 214
rect 938 204 950 206
rect 1005 184 1011 256
rect 1021 184 1027 236
rect 1117 184 1123 276
rect 1133 244 1139 276
rect 1229 264 1235 276
rect 804 177 812 183
rect 1204 177 1212 183
rect 772 157 780 163
rect 1053 144 1059 156
rect 1085 144 1091 156
rect 1261 144 1267 356
rect 1293 284 1299 296
rect 820 137 828 143
rect 1140 137 1148 143
rect 781 124 787 136
rect 861 124 867 136
rect 820 117 828 123
rect 212 97 220 103
rect 13 84 19 96
rect 346 14 358 16
rect 336 6 338 14
rect 346 6 348 14
rect 356 6 358 14
rect 366 6 368 14
rect 346 4 358 6
rect 541 -37 547 36
rect 541 -43 563 -37
rect 989 -43 995 116
rect 1053 24 1059 136
rect 1124 117 1132 123
rect 1149 24 1155 136
rect 1021 -43 1027 16
rect 1181 -43 1187 16
<< m3contact >>
rect 172 616 180 624
rect 156 576 164 584
rect 220 576 228 584
rect 316 616 324 624
rect 396 616 404 624
rect 396 596 404 604
rect 428 596 436 604
rect 444 556 452 564
rect 540 556 548 564
rect 636 556 644 564
rect 764 556 772 564
rect 796 556 804 564
rect 920 606 928 614
rect 930 606 938 614
rect 940 606 948 614
rect 950 606 958 614
rect 960 606 968 614
rect 972 556 980 564
rect 556 536 564 544
rect 588 536 596 544
rect 684 536 692 544
rect 828 536 836 544
rect 28 516 36 524
rect 924 516 932 524
rect 1036 516 1044 524
rect 1068 516 1076 524
rect 12 496 20 504
rect 60 496 68 504
rect 108 496 116 504
rect 380 436 388 444
rect 412 436 420 444
rect 328 406 336 414
rect 338 406 346 414
rect 348 406 356 414
rect 358 406 366 414
rect 368 406 376 414
rect 108 316 116 324
rect 156 296 164 304
rect 172 296 180 304
rect 268 296 276 304
rect 284 296 292 304
rect 364 296 372 304
rect 12 276 20 284
rect 124 276 132 284
rect 156 276 164 284
rect 332 276 340 284
rect 412 276 420 284
rect 12 256 20 264
rect 140 256 148 264
rect 188 256 196 264
rect 204 256 212 264
rect 268 256 276 264
rect 220 236 228 244
rect 172 156 180 164
rect 204 136 212 144
rect 284 176 292 184
rect 156 116 164 124
rect 492 436 500 444
rect 556 436 564 444
rect 444 336 452 344
rect 524 316 532 324
rect 716 496 724 504
rect 780 496 788 504
rect 828 496 836 504
rect 604 296 612 304
rect 1164 516 1172 524
rect 1068 376 1076 384
rect 1132 376 1140 384
rect 860 336 868 344
rect 908 336 916 344
rect 812 316 820 324
rect 844 316 852 324
rect 780 296 788 304
rect 860 296 868 304
rect 1180 356 1188 364
rect 1148 336 1156 344
rect 1196 316 1204 324
rect 668 276 676 284
rect 780 276 788 284
rect 908 276 916 284
rect 956 276 964 284
rect 1052 276 1060 284
rect 1292 496 1300 504
rect 1260 356 1268 364
rect 1244 316 1252 324
rect 1228 296 1236 304
rect 1116 276 1124 284
rect 460 256 468 264
rect 652 256 660 264
rect 780 256 788 264
rect 860 256 868 264
rect 1084 256 1092 264
rect 476 236 484 244
rect 732 236 740 244
rect 396 176 404 184
rect 428 176 436 184
rect 444 176 452 184
rect 588 176 596 184
rect 444 156 452 164
rect 460 136 468 144
rect 716 156 724 164
rect 924 236 932 244
rect 920 206 928 214
rect 930 206 938 214
rect 940 206 948 214
rect 950 206 958 214
rect 960 206 968 214
rect 1020 236 1028 244
rect 1228 256 1236 264
rect 1132 236 1140 244
rect 812 176 820 184
rect 1004 176 1012 184
rect 1212 176 1220 184
rect 780 156 788 164
rect 1052 156 1060 164
rect 1292 296 1300 304
rect 780 136 788 144
rect 812 136 820 144
rect 1084 136 1092 144
rect 1132 136 1140 144
rect 828 116 836 124
rect 860 116 868 124
rect 12 96 20 104
rect 220 96 228 104
rect 300 96 308 104
rect 328 6 336 14
rect 338 6 346 14
rect 348 6 356 14
rect 358 6 366 14
rect 368 6 376 14
rect 1116 116 1124 124
rect 1020 16 1028 24
rect 1052 16 1060 24
rect 1148 16 1156 24
rect 1180 16 1188 24
<< metal3 >>
rect 180 617 316 623
rect 324 617 396 623
rect 938 614 950 616
rect 938 604 950 606
rect 404 597 428 603
rect 164 577 220 583
rect 548 557 636 563
rect 772 557 796 563
rect 445 543 451 556
rect 445 537 556 543
rect 596 537 684 543
rect 973 543 979 556
rect 836 537 979 543
rect 36 517 115 523
rect 109 504 115 517
rect 932 517 1036 523
rect 1076 517 1164 523
rect -51 497 12 503
rect 68 497 76 503
rect 724 497 780 503
rect 788 497 828 503
rect 1300 497 1347 503
rect 388 437 412 443
rect 500 437 556 443
rect 346 414 358 416
rect 346 404 358 406
rect 1076 377 1132 383
rect 1188 357 1260 363
rect 1268 357 1347 363
rect 845 337 860 343
rect 868 337 908 343
rect 1140 337 1148 343
rect -51 317 108 323
rect 445 323 451 336
rect 445 317 524 323
rect 820 317 844 323
rect 1204 317 1244 323
rect 164 297 172 303
rect 180 297 268 303
rect 292 297 364 303
rect 596 297 604 303
rect 788 297 860 303
rect 1204 297 1228 303
rect 1300 297 1347 303
rect -51 277 12 283
rect 132 277 156 283
rect 340 277 412 283
rect 676 277 780 283
rect 916 277 956 283
rect 964 277 1052 283
rect 1124 277 1235 283
rect 1229 264 1235 277
rect 20 257 140 263
rect 196 257 204 263
rect 276 257 460 263
rect 660 257 780 263
rect 868 257 1084 263
rect 205 237 220 243
rect 228 237 476 243
rect 740 237 924 243
rect 1028 237 1132 243
rect 938 214 950 216
rect 938 204 950 206
rect 292 177 396 183
rect 436 177 444 183
rect 797 177 812 183
rect 820 177 1004 183
rect 1204 177 1212 183
rect 589 164 595 176
rect 68 157 172 163
rect 180 157 444 163
rect 765 157 780 163
rect 788 157 1052 163
rect 157 137 204 143
rect 157 124 163 137
rect 717 143 723 156
rect 468 137 723 143
rect 788 137 812 143
rect 1092 137 1132 143
rect 836 117 860 123
rect 1124 117 1132 123
rect -51 97 12 103
rect 228 97 300 103
rect 1028 17 1052 23
rect 1156 17 1180 23
rect 346 14 358 16
rect 346 4 358 6
<< m4contact >>
rect 922 606 928 614
rect 928 606 930 614
rect 934 606 938 614
rect 938 606 940 614
rect 940 606 942 614
rect 946 606 948 614
rect 948 606 950 614
rect 950 606 954 614
rect 958 606 960 614
rect 960 606 966 614
rect 76 496 84 504
rect 330 406 336 414
rect 336 406 338 414
rect 342 406 346 414
rect 346 406 348 414
rect 348 406 350 414
rect 354 406 356 414
rect 356 406 358 414
rect 358 406 362 414
rect 366 406 368 414
rect 368 406 374 414
rect 1132 336 1140 344
rect 588 296 596 304
rect 1196 296 1204 304
rect 922 206 928 214
rect 928 206 930 214
rect 934 206 938 214
rect 938 206 940 214
rect 940 206 942 214
rect 946 206 948 214
rect 948 206 950 214
rect 950 206 954 214
rect 958 206 960 214
rect 960 206 966 214
rect 1196 176 1204 184
rect 60 156 68 164
rect 588 156 596 164
rect 1132 116 1140 124
rect 330 6 336 14
rect 336 6 338 14
rect 342 6 346 14
rect 346 6 348 14
rect 348 6 350 14
rect 354 6 356 14
rect 356 6 358 14
rect 358 6 362 14
rect 366 6 368 14
rect 368 6 374 14
<< metal4 >>
rect 938 614 950 616
rect 938 604 950 606
rect 61 497 76 503
rect 61 164 67 497
rect 346 414 358 416
rect 346 404 358 406
rect 589 164 595 296
rect 938 214 950 216
rect 938 204 950 206
rect 1133 124 1139 336
rect 1197 184 1203 296
rect 346 14 358 16
rect 346 4 358 6
<< m5contact >>
rect 920 606 922 614
rect 922 606 928 614
rect 930 606 934 614
rect 934 606 938 614
rect 940 606 942 614
rect 942 606 946 614
rect 946 606 948 614
rect 950 606 954 614
rect 954 606 958 614
rect 960 606 966 614
rect 966 606 968 614
rect 328 406 330 414
rect 330 406 336 414
rect 338 406 342 414
rect 342 406 346 414
rect 348 406 350 414
rect 350 406 354 414
rect 354 406 356 414
rect 358 406 362 414
rect 362 406 366 414
rect 368 406 374 414
rect 374 406 376 414
rect 920 206 922 214
rect 922 206 928 214
rect 930 206 934 214
rect 934 206 938 214
rect 940 206 942 214
rect 942 206 946 214
rect 946 206 948 214
rect 950 206 954 214
rect 954 206 958 214
rect 960 206 966 214
rect 966 206 968 214
rect 328 6 330 14
rect 330 6 336 14
rect 338 6 342 14
rect 342 6 346 14
rect 348 6 350 14
rect 350 6 354 14
rect 354 6 356 14
rect 358 6 362 14
rect 362 6 366 14
rect 368 6 374 14
rect 374 6 376 14
<< metal5 >>
rect 938 615 950 616
rect 942 614 946 615
rect 928 606 930 614
rect 958 606 960 614
rect 942 605 946 606
rect 938 604 950 605
rect 346 415 358 416
rect 350 414 354 415
rect 336 406 338 414
rect 366 406 368 414
rect 350 405 354 406
rect 346 404 358 405
rect 938 215 950 216
rect 942 214 946 215
rect 928 206 930 214
rect 958 206 960 214
rect 942 205 946 206
rect 938 204 950 205
rect 346 15 358 16
rect 350 14 354 15
rect 336 6 338 14
rect 366 6 368 14
rect 350 5 354 6
rect 346 4 358 5
<< m6contact >>
rect 932 614 942 615
rect 946 614 956 615
rect 932 606 938 614
rect 938 606 940 614
rect 940 606 942 614
rect 946 606 948 614
rect 948 606 950 614
rect 950 606 956 614
rect 932 605 942 606
rect 946 605 956 606
rect 340 414 350 415
rect 354 414 364 415
rect 340 406 346 414
rect 346 406 348 414
rect 348 406 350 414
rect 354 406 356 414
rect 356 406 358 414
rect 358 406 364 414
rect 340 405 350 406
rect 354 405 364 406
rect 932 214 942 215
rect 946 214 956 215
rect 932 206 938 214
rect 938 206 940 214
rect 940 206 942 214
rect 946 206 948 214
rect 948 206 950 214
rect 950 206 956 214
rect 932 205 942 206
rect 946 205 956 206
rect 340 14 350 15
rect 354 14 364 15
rect 340 6 346 14
rect 346 6 348 14
rect 348 6 350 14
rect 354 6 356 14
rect 356 6 358 14
rect 358 6 364 14
rect 340 5 350 6
rect 354 5 364 6
<< metal6 >>
rect 328 415 376 615
rect 328 405 340 415
rect 350 405 354 415
rect 364 405 376 415
rect 328 15 376 405
rect 328 5 340 15
rect 350 5 354 15
rect 364 5 376 15
rect 328 -10 376 5
rect 920 605 932 615
rect 942 605 946 615
rect 956 605 968 615
rect 920 215 968 605
rect 920 205 932 215
rect 942 205 946 215
rect 956 205 968 215
rect 920 -10 968 205
use BUFX2  _31_
timestamp 1591289005
transform -1 0 56 0 -1 210
box -4 -6 52 206
use XOR2X1  _89_
timestamp 1591289005
transform -1 0 168 0 -1 210
box -4 -6 116 206
use XOR2X1  _61_
timestamp 1591289005
transform -1 0 120 0 1 210
box -4 -6 116 206
use INVX1  _58_
timestamp 1591289005
transform 1 0 120 0 1 210
box -4 -6 36 206
use NAND2X1  _76_
timestamp 1591289005
transform 1 0 168 0 -1 210
box -4 -6 52 206
use NAND2X1  _77_
timestamp 1591289005
transform -1 0 264 0 -1 210
box -4 -6 52 206
use INVX1  _57_
timestamp 1591289005
transform 1 0 152 0 1 210
box -4 -6 36 206
use NOR2X1  _59_
timestamp 1591289005
transform -1 0 232 0 1 210
box -4 -6 52 206
use NAND2X1  _60_
timestamp 1591289005
transform 1 0 232 0 1 210
box -4 -6 52 206
use INVX1  _75_
timestamp 1591289005
transform -1 0 296 0 -1 210
box -4 -6 36 206
use AND2X2  _81_
timestamp 1591289005
transform 1 0 296 0 -1 210
box -4 -6 68 206
use NAND2X1  _55_
timestamp 1591289005
transform -1 0 328 0 1 210
box -4 -6 52 206
use FILL  SFILL1800x50
timestamp 1591289005
transform -1 0 376 0 -1 210
box -4 -6 20 206
use FILL  SFILL1640x1050
timestamp 1591289005
transform 1 0 328 0 1 210
box -4 -6 20 206
use FILL  SFILL1720x1050
timestamp 1591289005
transform 1 0 344 0 1 210
box -4 -6 20 206
use FILL  SFILL1800x1050
timestamp 1591289005
transform 1 0 360 0 1 210
box -4 -6 20 206
use NAND2X1  _83_
timestamp 1591289005
transform -1 0 456 0 -1 210
box -4 -6 52 206
use NAND2X1  _84_
timestamp 1591289005
transform -1 0 504 0 -1 210
box -4 -6 52 206
use NOR2X1  _54_
timestamp 1591289005
transform -1 0 424 0 1 210
box -4 -6 52 206
use NAND2X1  _79_
timestamp 1591289005
transform 1 0 424 0 1 210
box -4 -6 52 206
use INVX1  _78_
timestamp 1591289005
transform 1 0 472 0 1 210
box -4 -6 36 206
use FILL  SFILL1880x50
timestamp 1591289005
transform -1 0 392 0 -1 210
box -4 -6 20 206
use FILL  SFILL1960x50
timestamp 1591289005
transform -1 0 408 0 -1 210
box -4 -6 20 206
use INVX1  _82_
timestamp 1591289005
transform -1 0 536 0 -1 210
box -4 -6 36 206
use BUFX2  _29_
timestamp 1591289005
transform -1 0 584 0 -1 210
box -4 -6 52 206
use INVX1  _68_
timestamp 1591289005
transform 1 0 584 0 -1 210
box -4 -6 36 206
use NAND2X1  _80_
timestamp 1591289005
transform 1 0 504 0 1 210
box -4 -6 52 206
use XOR2X1  _87_
timestamp 1591289005
transform -1 0 664 0 1 210
box -4 -6 116 206
use NAND2X1  _70_
timestamp 1591289005
transform 1 0 616 0 -1 210
box -4 -6 52 206
use INVX1  _72_
timestamp 1591289005
transform 1 0 664 0 -1 210
box -4 -6 36 206
use NAND2X1  _74_
timestamp 1591289005
transform 1 0 696 0 -1 210
box -4 -6 52 206
use NAND2X1  _69_
timestamp 1591289005
transform -1 0 712 0 1 210
box -4 -6 52 206
use INVX1  _65_
timestamp 1591289005
transform 1 0 712 0 1 210
box -4 -6 36 206
use INVX1  _37_
timestamp 1591289005
transform -1 0 776 0 -1 210
box -4 -6 36 206
use NOR2X1  _39_
timestamp 1591289005
transform 1 0 776 0 -1 210
box -4 -6 52 206
use NAND2X1  _40_
timestamp 1591289005
transform 1 0 824 0 -1 210
box -4 -6 52 206
use NAND2X1  _67_
timestamp 1591289005
transform 1 0 744 0 1 210
box -4 -6 52 206
use AND2X2  _71_
timestamp 1591289005
transform 1 0 792 0 1 210
box -4 -6 68 206
use INVX1  _38_
timestamp 1591289005
transform -1 0 904 0 -1 210
box -4 -6 36 206
use XOR2X1  _41_
timestamp 1591289005
transform -1 0 1064 0 -1 210
box -4 -6 116 206
use NAND2X1  _66_
timestamp 1591289005
transform -1 0 904 0 1 210
box -4 -6 52 206
use NAND2X1  _73_
timestamp 1591289005
transform -1 0 952 0 1 210
box -4 -6 52 206
use FILL  SFILL4520x50
timestamp 1591289005
transform -1 0 920 0 -1 210
box -4 -6 20 206
use FILL  SFILL4600x50
timestamp 1591289005
transform -1 0 936 0 -1 210
box -4 -6 20 206
use FILL  SFILL4680x50
timestamp 1591289005
transform -1 0 952 0 -1 210
box -4 -6 20 206
use FILL  SFILL4760x1050
timestamp 1591289005
transform 1 0 952 0 1 210
box -4 -6 20 206
use FILL  SFILL4840x1050
timestamp 1591289005
transform 1 0 968 0 1 210
box -4 -6 20 206
use INVX1  _33_
timestamp 1591289005
transform -1 0 1096 0 -1 210
box -4 -6 36 206
use INVX1  _62_
timestamp 1591289005
transform 1 0 1000 0 1 210
box -4 -6 36 206
use NAND2X1  _64_
timestamp 1591289005
transform 1 0 1032 0 1 210
box -4 -6 52 206
use NAND2X1  _63_
timestamp 1591289005
transform -1 0 1128 0 1 210
box -4 -6 52 206
use FILL  SFILL4920x1050
timestamp 1591289005
transform 1 0 984 0 1 210
box -4 -6 20 206
use NOR2X1  _35_
timestamp 1591289005
transform 1 0 1096 0 -1 210
box -4 -6 52 206
use XOR2X1  _36_
timestamp 1591289005
transform 1 0 1144 0 -1 210
box -4 -6 116 206
use XOR2X1  _85_
timestamp 1591289005
transform -1 0 1240 0 1 210
box -4 -6 116 206
use BUFX2  _27_
timestamp 1591289005
transform 1 0 1240 0 1 210
box -4 -6 52 206
use FILL  FILL5800x50
timestamp 1591289005
transform -1 0 1272 0 -1 210
box -4 -6 20 206
use FILL  FILL5880x50
timestamp 1591289005
transform -1 0 1288 0 -1 210
box -4 -6 20 206
use BUFX2  _30_
timestamp 1591289005
transform -1 0 56 0 -1 610
box -4 -6 52 206
use XOR2X1  _88_
timestamp 1591289005
transform 1 0 56 0 -1 610
box -4 -6 116 206
use XOR2X1  _56_
timestamp 1591289005
transform 1 0 168 0 -1 610
box -4 -6 116 206
use INVX1  _53_
timestamp 1591289005
transform 1 0 280 0 -1 610
box -4 -6 36 206
use INVX1  _52_
timestamp 1591289005
transform 1 0 312 0 -1 610
box -4 -6 36 206
use FILL  SFILL1720x2050
timestamp 1591289005
transform -1 0 360 0 -1 610
box -4 -6 20 206
use FILL  SFILL1800x2050
timestamp 1591289005
transform -1 0 376 0 -1 610
box -4 -6 20 206
use BUFX2  _32_
timestamp 1591289005
transform -1 0 440 0 -1 610
box -4 -6 52 206
use XOR2X1  _51_
timestamp 1591289005
transform 1 0 440 0 -1 610
box -4 -6 116 206
use FILL  SFILL1880x2050
timestamp 1591289005
transform -1 0 392 0 -1 610
box -4 -6 20 206
use INVX1  _47_
timestamp 1591289005
transform 1 0 552 0 -1 610
box -4 -6 36 206
use NOR2X1  _49_
timestamp 1591289005
transform 1 0 584 0 -1 610
box -4 -6 52 206
use INVX1  _48_
timestamp 1591289005
transform 1 0 632 0 -1 610
box -4 -6 36 206
use NAND2X1  _50_
timestamp 1591289005
transform -1 0 712 0 -1 610
box -4 -6 52 206
use NOR2X1  _44_
timestamp 1591289005
transform -1 0 760 0 -1 610
box -4 -6 52 206
use NAND2X1  _45_
timestamp 1591289005
transform -1 0 808 0 -1 610
box -4 -6 52 206
use INVX1  _42_
timestamp 1591289005
transform -1 0 840 0 -1 610
box -4 -6 36 206
use INVX1  _43_
timestamp 1591289005
transform -1 0 872 0 -1 610
box -4 -6 36 206
use XOR2X1  _46_
timestamp 1591289005
transform -1 0 984 0 -1 610
box -4 -6 116 206
use XOR2X1  _86_
timestamp 1591289005
transform -1 0 1144 0 -1 610
box -4 -6 116 206
use FILL  SFILL4920x2050
timestamp 1591289005
transform -1 0 1000 0 -1 610
box -4 -6 20 206
use FILL  SFILL5000x2050
timestamp 1591289005
transform -1 0 1016 0 -1 610
box -4 -6 20 206
use FILL  SFILL5080x2050
timestamp 1591289005
transform -1 0 1032 0 -1 610
box -4 -6 20 206
use INVX1  _34_
timestamp 1591289005
transform -1 0 1176 0 -1 610
box -4 -6 36 206
use BUFX2  _28_
timestamp 1591289005
transform 1 0 1176 0 -1 610
box -4 -6 52 206
use BUFX2  _26_
timestamp 1591289005
transform 1 0 1224 0 -1 610
box -4 -6 52 206
use FILL  FILL5880x2050
timestamp 1591289005
transform -1 0 1288 0 -1 610
box -4 -6 20 206
<< labels >>
flabel metal6 s 920 -10 968 0 7 FreeSans 48 270 0 0 gnd
port 0 nsew
flabel metal6 s 328 -10 376 0 7 FreeSans 48 270 0 0 vdd
port 1 nsew
flabel metal2 s 429 677 435 683 3 FreeSans 48 90 0 0 s[6]
port 2 nsew
flabel metal3 s -51 97 -45 103 7 FreeSans 48 0 0 0 s[5]
port 3 nsew
flabel metal3 s -51 497 -45 503 7 FreeSans 48 0 0 0 s[4]
port 4 nsew
flabel metal2 s 557 -43 563 -37 7 FreeSans 48 270 0 0 s[3]
port 5 nsew
flabel metal2 s 1197 677 1203 683 3 FreeSans 48 90 0 0 s[2]
port 6 nsew
flabel metal3 s 1341 297 1347 303 3 FreeSans 48 0 0 0 s[1]
port 7 nsew
flabel metal3 s 1341 497 1347 503 3 FreeSans 48 0 0 0 s[0]
port 8 nsew
flabel metal3 s -51 277 -45 283 7 FreeSans 48 0 0 0 x[5]
port 9 nsew
flabel metal2 s 285 677 291 683 3 FreeSans 48 90 0 0 x[4]
port 10 nsew
flabel metal2 s 637 677 643 683 3 FreeSans 48 90 0 0 x[3]
port 11 nsew
flabel metal2 s 877 677 883 683 3 FreeSans 48 90 0 0 x[2]
port 12 nsew
flabel metal2 s 989 -43 995 -37 7 FreeSans 48 270 0 0 x[1]
port 13 nsew
flabel metal3 s 1341 357 1347 363 3 FreeSans 48 0 0 0 x[0]
port 14 nsew
flabel metal3 s -51 317 -45 323 7 FreeSans 48 0 0 0 y[5]
port 15 nsew
flabel metal2 s 397 677 403 683 3 FreeSans 48 90 0 0 y[4]
port 16 nsew
flabel metal2 s 557 677 563 683 3 FreeSans 48 90 0 0 y[3]
port 17 nsew
flabel metal2 s 829 677 835 683 3 FreeSans 48 90 0 0 y[2]
port 18 nsew
flabel metal2 s 1021 -43 1027 -37 7 FreeSans 48 270 0 0 y[1]
port 19 nsew
flabel metal2 s 1181 -43 1187 -37 7 FreeSans 48 270 0 0 y[0]
port 20 nsew
<< end >>
