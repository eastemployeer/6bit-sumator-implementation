VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 1000 ;
END UNITS

MACRO single_generate
  CLASS BLOCK ;
  FOREIGN single_generate ;
  ORIGIN 2.600000 0.600000 ;
  SIZE 31.600000 BY 14.800000 ;
  PIN gnd
    USE GROUND ;
    PORT
      LAYER metal1 ;
        RECT 0.200000 10.200000 26.200001 10.800000 ;
        RECT 1.400000 7.900000 1.800000 10.200000 ;
        RECT 3.900000 9.900001 4.300000 10.200000 ;
        RECT 3.800000 8.200000 4.300000 9.900001 ;
        RECT 6.900000 8.200000 7.400000 10.200000 ;
        RECT 11.000000 8.900001 11.400001 10.200000 ;
        RECT 13.400001 7.900000 13.800000 10.200000 ;
        RECT 15.000000 8.900001 15.400001 10.200000 ;
        RECT 16.600000 8.900001 17.000000 10.200000 ;
        RECT 18.200001 8.900001 18.600000 10.200000 ;
        RECT 21.400000 7.900000 21.800001 10.200000 ;
        RECT 24.600000 7.900000 25.000000 10.200000 ;
      LAYER via1 ;
        RECT 17.200001 10.300000 17.600000 10.700000 ;
        RECT 17.700001 10.300000 18.100000 10.700000 ;
        RECT 18.200001 10.300000 18.600000 10.700000 ;
        RECT 18.700001 10.300000 19.100000 10.700000 ;
        RECT 19.200001 10.300000 19.600000 10.700000 ;
      LAYER metal2 ;
        RECT 18.100000 10.700000 18.700001 10.800000 ;
        RECT 17.200001 10.300000 19.600000 10.700000 ;
        RECT 18.100000 10.200000 18.700001 10.300000 ;
      LAYER via2 ;
        RECT 17.700001 10.300000 18.100000 10.700000 ;
        RECT 18.200001 10.300000 18.600000 10.700000 ;
        RECT 18.700001 10.300000 19.100000 10.700000 ;
        RECT 19.200001 10.300000 19.600000 10.700000 ;
      LAYER metal3 ;
        RECT 18.100000 10.700000 18.700001 10.800000 ;
        RECT 17.200001 10.300000 19.600000 10.700000 ;
        RECT 18.100000 10.200000 18.700001 10.300000 ;
      LAYER via3 ;
        RECT 17.300001 10.300000 17.700001 10.700000 ;
        RECT 17.900000 10.300000 18.300001 10.700000 ;
        RECT 18.500000 10.300000 18.900000 10.700000 ;
        RECT 19.100000 10.300000 19.500000 10.700000 ;
      LAYER metal4 ;
        RECT 18.100000 10.700000 18.700001 10.800000 ;
        RECT 17.200001 10.300000 19.600000 10.700000 ;
        RECT 18.100000 10.200000 18.700001 10.300000 ;
      LAYER via4 ;
        RECT 17.200001 10.300000 17.600000 10.700000 ;
        RECT 17.700001 10.300000 18.100000 10.700000 ;
        RECT 18.200001 10.300000 18.600000 10.700000 ;
        RECT 18.700001 10.300000 19.100000 10.700000 ;
        RECT 19.200001 10.300000 19.600000 10.700000 ;
      LAYER metal5 ;
        RECT 18.100000 10.700000 18.700001 10.800000 ;
        RECT 17.200001 10.300000 19.600000 10.700000 ;
        RECT 17.800001 10.200000 19.000000 10.300000 ;
      LAYER via5 ;
        RECT 18.500000 10.200000 19.000000 10.700000 ;
      LAYER metal6 ;
        RECT 17.200001 -0.600000 19.600000 10.700000 ;
    END
  END gnd
  PIN vdd
    USE POWER ;
    PORT
      LAYER metal1 ;
        RECT 1.400000 0.800000 1.800000 4.500000 ;
        RECT 3.800000 1.100000 4.300000 4.400000 ;
        RECT 3.900000 0.800000 4.300000 1.100000 ;
        RECT 6.900000 0.800000 7.400000 4.400000 ;
        RECT 11.000000 0.800000 11.400001 3.100000 ;
        RECT 13.400001 0.800000 13.800000 4.500000 ;
        RECT 15.000000 0.800000 15.400001 3.100000 ;
        RECT 16.600000 0.800000 17.000000 5.100000 ;
        RECT 21.400000 0.800000 21.800001 3.100000 ;
        RECT 23.000000 0.800000 23.400000 3.100000 ;
        RECT 24.600000 0.800000 25.000000 4.500000 ;
        RECT 0.200000 0.200000 26.200001 0.800000 ;
      LAYER via1 ;
        RECT 6.800000 0.300000 7.200000 0.700000 ;
        RECT 7.300000 0.300000 7.700000 0.700000 ;
        RECT 7.800000 0.300000 8.200000 0.700000 ;
        RECT 8.300000 0.300000 8.700000 0.700000 ;
        RECT 8.800000 0.300000 9.200000 0.700000 ;
      LAYER metal2 ;
        RECT 7.700000 0.700000 8.300000 0.800000 ;
        RECT 6.800000 0.300000 9.200000 0.700000 ;
        RECT 7.700000 0.200000 8.300000 0.300000 ;
      LAYER via2 ;
        RECT 7.300000 0.300000 7.700000 0.700000 ;
        RECT 7.800000 0.300000 8.200000 0.700000 ;
        RECT 8.300000 0.300000 8.700000 0.700000 ;
        RECT 8.800000 0.300000 9.200000 0.700000 ;
      LAYER metal3 ;
        RECT 7.700000 0.700000 8.300000 0.800000 ;
        RECT 6.800000 0.300000 9.200000 0.700000 ;
        RECT 7.700000 0.200000 8.300000 0.300000 ;
      LAYER via3 ;
        RECT 6.900000 0.300000 7.300000 0.700000 ;
        RECT 7.500000 0.300000 7.900000 0.700000 ;
        RECT 8.100000 0.300000 8.500000 0.700000 ;
        RECT 8.700000 0.300000 9.100000 0.700000 ;
      LAYER metal4 ;
        RECT 7.700000 0.700000 8.300000 0.800000 ;
        RECT 6.800000 0.300000 9.200000 0.700000 ;
        RECT 7.700000 0.200000 8.300000 0.300000 ;
      LAYER via4 ;
        RECT 6.800000 0.300000 7.200000 0.700000 ;
        RECT 7.300000 0.300000 7.700000 0.700000 ;
        RECT 7.800000 0.300000 8.200000 0.700000 ;
        RECT 8.300000 0.300000 8.700000 0.700000 ;
        RECT 8.800000 0.300000 9.200000 0.700000 ;
      LAYER metal5 ;
        RECT 7.700000 0.700000 8.300000 0.800000 ;
        RECT 6.800000 0.300000 9.200000 0.700000 ;
        RECT 7.400000 0.200000 8.600000 0.300000 ;
      LAYER via5 ;
        RECT 8.100000 0.200000 8.600000 0.700000 ;
      LAYER metal6 ;
        RECT 6.800000 -0.600000 9.200000 10.700000 ;
    END
  END vdd
  PIN g
    PORT
      LAYER metal1 ;
        RECT 12.600000 6.200000 13.000000 9.900001 ;
        RECT 12.600000 5.100000 12.900001 6.200000 ;
        RECT 12.600000 1.100000 13.000000 5.100000 ;
      LAYER via1 ;
        RECT 12.600000 8.800000 13.000000 9.200000 ;
      LAYER metal2 ;
        RECT 13.400001 14.100000 13.800000 14.200000 ;
        RECT 12.600000 13.800000 13.800000 14.100000 ;
        RECT 12.600000 9.200000 12.900001 13.800000 ;
        RECT 12.600000 8.800000 13.000000 9.200000 ;
    END
  END g
  PIN h
    PORT
      LAYER metal1 ;
        RECT 0.600000 6.200000 1.000000 9.900001 ;
        RECT 0.600000 5.100000 0.900000 6.200000 ;
        RECT 0.600000 1.100000 1.000000 5.100000 ;
      LAYER via1 ;
        RECT 0.600000 3.800000 1.000000 4.200000 ;
      LAYER metal2 ;
        RECT 0.600000 4.800000 1.000000 5.200000 ;
        RECT 0.600000 4.200000 0.900000 4.800000 ;
        RECT 0.600000 3.800000 1.000000 4.200000 ;
      LAYER metal3 ;
        RECT -2.600000 5.100000 -2.200000 5.200000 ;
        RECT 0.600000 5.100000 1.000000 5.200000 ;
        RECT -2.600000 4.800000 1.000000 5.100000 ;
    END
  END h
  PIN p
    PORT
      LAYER metal1 ;
        RECT 25.400000 6.200000 25.800001 9.900001 ;
        RECT 25.500000 5.100000 25.800001 6.200000 ;
        RECT 25.400000 4.100000 25.800001 5.100000 ;
        RECT 26.200001 4.100000 26.600000 4.200000 ;
        RECT 25.400000 3.800000 26.600000 4.100000 ;
        RECT 25.400000 1.100000 25.800001 3.800000 ;
      LAYER via1 ;
        RECT 26.200001 3.800000 26.600000 4.200000 ;
      LAYER metal2 ;
        RECT 26.200001 4.800000 26.600000 5.200000 ;
        RECT 26.200001 4.200000 26.500000 4.800000 ;
        RECT 26.200001 3.800000 26.600000 4.200000 ;
      LAYER metal3 ;
        RECT 26.200001 5.100000 26.600000 5.200000 ;
        RECT 28.600000 5.100000 29.000000 5.200000 ;
        RECT 26.200001 4.800000 29.000000 5.100000 ;
    END
  END p
  PIN x
    PORT
      LAYER metal1 ;
        RECT 10.200000 8.100000 10.600000 8.200000 ;
        RECT 11.000000 8.100000 11.400001 8.600000 ;
        RECT 10.200000 7.800000 11.400001 8.100000 ;
        RECT 7.400000 7.100000 8.200000 7.200000 ;
        RECT 10.200000 7.100000 10.500000 7.800000 ;
        RECT 7.400000 6.800000 10.500000 7.100000 ;
      LAYER metal2 ;
        RECT 10.200000 13.800000 10.600000 14.200000 ;
        RECT 10.200000 8.200000 10.500000 13.800000 ;
        RECT 10.200000 7.800000 10.600000 8.200000 ;
    END
  END x
  PIN y
    PORT
      LAYER metal1 ;
        RECT 15.000000 7.800000 15.400001 8.600000 ;
        RECT 3.000000 7.100000 3.800000 7.200000 ;
        RECT 3.000000 7.000000 4.100000 7.100000 ;
        RECT 3.000000 6.800000 5.200000 7.000000 ;
        RECT 3.800000 6.700000 5.200000 6.800000 ;
        RECT 4.800000 6.600000 5.200000 6.700000 ;
      LAYER metal2 ;
        RECT 15.000000 13.800000 15.400001 14.200000 ;
        RECT 15.000000 8.200000 15.300000 13.800000 ;
        RECT 3.000000 7.800000 3.400000 8.200000 ;
        RECT 15.000000 7.800000 15.400001 8.200000 ;
        RECT 3.000000 7.200000 3.300000 7.800000 ;
        RECT 3.000000 6.800000 3.400000 7.200000 ;
      LAYER metal3 ;
        RECT 3.000000 8.100000 3.400000 8.200000 ;
        RECT 15.000000 8.100000 15.400001 8.200000 ;
        RECT 3.000000 7.800000 15.400001 8.100000 ;
    END
  END y
  OBS
      LAYER metal1 ;
        RECT 2.200000 7.600000 2.600000 9.900001 ;
        RECT 3.000000 7.900000 3.400000 9.900001 ;
        RECT 5.200000 8.100000 6.000000 9.900001 ;
        RECT 3.000000 7.600000 4.300000 7.900000 ;
        RECT 1.500000 7.300000 2.600000 7.600000 ;
        RECT 3.900000 7.500000 4.300000 7.600000 ;
        RECT 4.600000 7.400000 5.400000 7.800000 ;
        RECT 1.500000 5.800000 1.800000 7.300000 ;
        RECT 5.700000 7.100000 6.000000 8.100000 ;
        RECT 7.800000 7.900000 8.200000 9.900001 ;
        RECT 6.300000 7.400000 6.700000 7.800000 ;
        RECT 7.000000 7.600000 8.200000 7.900000 ;
        RECT 7.000000 7.500000 7.400000 7.600000 ;
        RECT 5.500000 6.800000 6.000000 7.100000 ;
        RECT 6.400000 7.200000 6.700000 7.400000 ;
        RECT 6.400000 6.800000 6.800000 7.200000 ;
        RECT 2.200000 6.100000 2.600000 6.600000 ;
        RECT 5.500000 6.200000 5.800000 6.800000 ;
        RECT 3.000000 6.100000 3.400000 6.200000 ;
        RECT 2.200000 5.800000 3.400000 6.100000 ;
        RECT 4.100000 6.100000 4.500000 6.200000 ;
        RECT 4.100000 5.800000 4.900000 6.100000 ;
        RECT 5.400000 5.800000 5.800000 6.200000 ;
        RECT 11.000000 6.100000 11.400001 6.200000 ;
        RECT 11.800000 6.100000 12.200000 9.900001 ;
        RECT 14.200000 7.600000 14.600000 9.900001 ;
        RECT 11.000000 5.800000 12.200000 6.100000 ;
        RECT 13.500000 7.300000 14.600000 7.600000 ;
        RECT 15.800000 8.100000 16.200001 9.900001 ;
        RECT 17.400000 8.900001 17.800001 9.900001 ;
        RECT 16.600000 8.100000 17.000000 8.600000 ;
        RECT 17.500000 8.200000 17.800001 8.900001 ;
        RECT 22.700001 8.200000 23.100000 9.900001 ;
        RECT 15.800000 7.800000 17.000000 8.100000 ;
        RECT 17.400000 7.800000 17.800001 8.200000 ;
        RECT 13.500000 5.800000 13.800000 7.300000 ;
        RECT 15.800000 7.100000 16.200001 7.800000 ;
        RECT 17.500000 7.200000 17.800001 7.800000 ;
        RECT 22.200001 7.900000 23.100000 8.200000 ;
        RECT 15.800000 6.800000 16.900000 7.100000 ;
        RECT 17.400000 6.800000 17.800001 7.200000 ;
        RECT 21.400000 6.800000 21.800001 7.600000 ;
        RECT 14.200000 6.100000 14.600000 6.600000 ;
        RECT 15.000000 6.100000 15.400001 6.200000 ;
        RECT 14.200000 5.800000 15.400001 6.100000 ;
        RECT 1.200000 5.400000 1.800000 5.800000 ;
        RECT 4.500000 5.700000 4.900000 5.800000 ;
        RECT 1.500000 5.100000 1.800000 5.400000 ;
        RECT 5.500000 5.100000 5.800000 5.800000 ;
        RECT 1.500000 4.800000 2.600000 5.100000 ;
        RECT 2.200000 1.100000 2.600000 4.800000 ;
        RECT 3.000000 4.800000 4.300000 5.100000 ;
        RECT 3.000000 1.100000 3.400000 4.800000 ;
        RECT 3.900000 4.700000 4.300000 4.800000 ;
        RECT 5.200000 1.100000 6.000000 5.100000 ;
        RECT 7.000000 4.800000 8.200000 5.100000 ;
        RECT 7.000000 4.700000 7.400000 4.800000 ;
        RECT 7.800000 1.100000 8.200000 4.800000 ;
        RECT 11.800000 1.100000 12.200000 5.800000 ;
        RECT 13.200000 5.400000 13.800000 5.800000 ;
        RECT 13.500000 5.100000 13.800000 5.400000 ;
        RECT 13.500000 4.800000 14.600000 5.100000 ;
        RECT 14.200000 1.100000 14.600000 4.800000 ;
        RECT 15.800000 1.100000 16.200001 6.800000 ;
        RECT 16.600000 6.200000 16.900000 6.800000 ;
        RECT 16.600000 5.800000 17.000000 6.200000 ;
        RECT 17.500000 5.100000 17.800001 6.800000 ;
        RECT 18.200001 5.400000 18.600000 6.200000 ;
        RECT 22.200001 6.100000 22.600000 7.900000 ;
        RECT 23.800001 7.600000 24.200001 9.900001 ;
        RECT 23.800001 7.300000 24.900000 7.600000 ;
        RECT 23.800001 6.100000 24.200001 6.600000 ;
        RECT 22.200001 5.800000 24.200001 6.100000 ;
        RECT 24.600000 5.800000 24.900000 7.300000 ;
        RECT 17.400000 4.700000 18.300001 5.100000 ;
        RECT 17.900000 1.100000 18.300001 4.700000 ;
        RECT 22.200001 1.100000 22.600000 5.800000 ;
        RECT 24.600000 5.400000 25.200001 5.800000 ;
        RECT 23.000000 4.400000 23.400000 5.200000 ;
        RECT 24.600000 5.100000 24.900000 5.400000 ;
        RECT 23.800001 4.800000 24.900000 5.100000 ;
        RECT 23.800001 1.100000 24.200001 4.800000 ;
      LAYER via1 ;
        RECT 3.000000 5.800000 3.400000 6.200000 ;
        RECT 15.000000 5.800000 15.400001 6.200000 ;
        RECT 18.200001 5.800000 18.600000 6.200000 ;
        RECT 23.000000 4.800000 23.400000 5.200000 ;
      LAYER metal2 ;
        RECT 16.600000 8.100000 17.000000 8.200000 ;
        RECT 17.400000 8.100000 17.800001 8.200000 ;
        RECT 3.900000 7.800000 4.300000 7.900000 ;
        RECT 3.900000 7.500000 6.700000 7.800000 ;
        RECT 7.000000 7.500000 7.400000 7.900000 ;
        RECT 16.600000 7.800000 17.800001 8.100000 ;
        RECT 2.200000 6.100000 2.600000 6.200000 ;
        RECT 3.000000 6.100000 3.400000 6.200000 ;
        RECT 2.200000 5.800000 3.400000 6.100000 ;
        RECT 3.900000 5.100000 4.200000 7.500000 ;
        RECT 4.600000 7.400000 5.000000 7.500000 ;
        RECT 6.300000 7.400000 6.700000 7.500000 ;
        RECT 7.100000 7.100000 7.400000 7.500000 ;
        RECT 4.600000 6.800000 7.400000 7.100000 ;
        RECT 4.600000 6.100000 4.900000 6.800000 ;
        RECT 4.500000 5.700000 4.900000 6.100000 ;
        RECT 5.400000 5.800000 5.800000 6.200000 ;
        RECT 5.400000 5.200000 5.700000 5.800000 ;
        RECT 3.900000 4.700000 4.300000 5.100000 ;
        RECT 5.400000 4.800000 5.800000 5.200000 ;
        RECT 7.100000 5.100000 7.400000 6.800000 ;
        RECT 15.000000 6.800000 15.400001 7.200000 ;
        RECT 16.600000 6.800000 17.000000 7.200000 ;
        RECT 20.600000 7.100000 21.000000 7.200000 ;
        RECT 21.400000 7.100000 21.800001 7.200000 ;
        RECT 20.600000 6.800000 21.800001 7.100000 ;
        RECT 15.000000 6.200000 15.300000 6.800000 ;
        RECT 16.600000 6.200000 16.900000 6.800000 ;
        RECT 11.000000 6.100000 11.400001 6.200000 ;
        RECT 11.800000 6.100000 12.200000 6.200000 ;
        RECT 11.000000 5.800000 12.200000 6.100000 ;
        RECT 15.000000 5.800000 15.400001 6.200000 ;
        RECT 16.600000 5.800000 17.000000 6.200000 ;
        RECT 17.400000 6.100000 17.800001 6.200000 ;
        RECT 18.200001 6.100000 18.600000 6.200000 ;
        RECT 17.400000 5.800000 18.600000 6.100000 ;
        RECT 23.000000 5.800000 23.400000 6.200000 ;
        RECT 7.000000 4.700000 7.400000 5.100000 ;
        RECT 23.000000 5.200000 23.300001 5.800000 ;
        RECT 23.000000 4.800000 23.400000 5.200000 ;
      LAYER via2 ;
        RECT 11.800000 5.800000 12.200000 6.200000 ;
      LAYER metal3 ;
        RECT 16.600000 8.100000 17.000000 8.200000 ;
        RECT 15.800000 7.800000 17.000000 8.100000 ;
        RECT 15.000000 7.100000 15.400001 7.200000 ;
        RECT 15.800000 7.100000 16.100000 7.800000 ;
        RECT 15.000000 6.800000 16.100000 7.100000 ;
        RECT 16.600000 7.100000 17.000000 7.200000 ;
        RECT 20.600000 7.100000 21.000000 7.200000 ;
        RECT 16.600000 6.800000 21.000000 7.100000 ;
        RECT 2.200000 6.100000 2.600000 6.200000 ;
        RECT 11.800000 6.100000 12.200000 6.200000 ;
        RECT 17.400000 6.100000 17.800001 6.200000 ;
        RECT 23.000000 6.100000 23.400000 6.200000 ;
        RECT 2.200000 5.800000 5.700000 6.100000 ;
        RECT 11.800000 5.800000 23.400000 6.100000 ;
        RECT 5.400000 5.200000 5.700000 5.800000 ;
        RECT 5.400000 4.800000 5.800000 5.200000 ;
  END
END single_generate
