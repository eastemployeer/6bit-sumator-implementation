VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 1000 ;
END UNITS

MACRO adder
  CLASS BLOCK ;
  FOREIGN adder ;
  ORIGIN 2.600000 2.200000 ;
  SIZE 70.000000 BY 36.400002 ;
  PIN gnd
    USE GROUND ;
    PORT
      LAYER metal1 ;
        RECT 0.200000 30.200001 64.599998 30.800001 ;
        RECT 1.400000 27.900000 1.800000 30.200001 ;
        RECT 3.900000 29.900000 4.300000 30.200001 ;
        RECT 3.800000 28.200001 4.300000 29.900000 ;
        RECT 6.900000 28.200001 7.400000 30.200001 ;
        RECT 9.500000 29.900000 9.900001 30.200001 ;
        RECT 9.400001 28.200001 9.900001 29.900000 ;
        RECT 12.500000 28.200001 13.000000 30.200001 ;
        RECT 14.200000 28.900000 14.600000 30.200001 ;
        RECT 15.800000 28.900000 16.200001 30.200001 ;
        RECT 20.600000 27.900000 21.000000 30.200001 ;
        RECT 23.100000 29.900000 23.500000 30.200001 ;
        RECT 23.000000 28.200001 23.500000 29.900000 ;
        RECT 26.100000 28.200001 26.600000 30.200001 ;
        RECT 27.800001 28.900000 28.200001 30.200001 ;
        RECT 29.400000 28.900000 29.800001 30.200001 ;
        RECT 31.000000 28.900000 31.400000 30.200001 ;
        RECT 31.800001 28.900000 32.200001 30.200001 ;
        RECT 35.000000 27.900000 35.400002 30.200001 ;
        RECT 35.799999 28.900000 36.200001 30.200001 ;
        RECT 37.400002 28.900000 37.799999 30.200001 ;
        RECT 39.799999 27.900000 40.200001 30.200001 ;
        RECT 41.400002 28.900000 41.799999 30.200001 ;
        RECT 43.000000 28.900000 43.400002 30.200001 ;
        RECT 44.600002 28.200001 45.100002 30.200001 ;
        RECT 47.700001 29.900000 48.100002 30.200001 ;
        RECT 47.700001 28.200001 48.200001 29.900000 ;
        RECT 52.600002 28.200001 53.100002 30.200001 ;
        RECT 55.700001 29.900000 56.100002 30.200001 ;
        RECT 55.700001 28.200001 56.200001 29.900000 ;
        RECT 58.200001 28.900000 58.600002 30.200001 ;
        RECT 59.799999 27.900000 60.200001 30.200001 ;
        RECT 62.200001 27.900000 62.600002 30.200001 ;
        RECT 1.400000 10.800000 1.900000 12.800000 ;
        RECT 4.500000 11.100000 5.000000 12.800000 ;
        RECT 4.500000 10.800000 4.900000 11.100000 ;
        RECT 6.200000 10.800000 6.600000 12.100000 ;
        RECT 7.800000 10.800000 8.200000 12.100000 ;
        RECT 9.400001 10.800000 9.800000 12.100000 ;
        RECT 11.000000 10.800000 11.400001 12.100000 ;
        RECT 11.800000 10.800000 12.200000 13.100000 ;
        RECT 15.800000 10.800000 16.200001 13.100000 ;
        RECT 19.000000 10.800000 19.400000 12.100000 ;
        RECT 20.600000 10.800000 21.000000 12.100000 ;
        RECT 21.400000 10.800000 21.800001 13.100000 ;
        RECT 23.800001 10.800000 24.200001 12.100000 ;
        RECT 25.400000 10.800000 25.800001 13.100000 ;
        RECT 28.600000 10.800000 29.100000 12.800000 ;
        RECT 31.700001 11.100000 32.200001 12.800000 ;
        RECT 31.700001 10.800000 32.100002 11.100000 ;
        RECT 35.000000 10.800000 35.400002 13.100000 ;
        RECT 35.799999 10.800000 36.200001 12.100000 ;
        RECT 37.400002 10.800000 37.799999 13.100000 ;
        RECT 41.100002 10.800000 41.500000 13.000000 ;
        RECT 44.600002 10.800000 45.000000 13.100000 ;
        RECT 47.000000 10.800000 47.400002 13.100000 ;
        RECT 50.200001 10.800000 50.600002 12.100000 ;
        RECT 51.799999 10.800000 52.200001 13.100000 ;
        RECT 55.799999 10.800000 56.200001 13.100000 ;
        RECT 57.400002 10.800000 57.900002 12.800000 ;
        RECT 60.500000 11.100000 61.000000 12.800000 ;
        RECT 60.500000 10.800000 60.900002 11.100000 ;
        RECT 63.000000 10.800000 63.400002 13.100000 ;
        RECT 0.200000 10.200000 64.599998 10.800000 ;
        RECT 1.400000 7.900000 1.800000 10.200000 ;
        RECT 3.800000 8.200000 4.300000 10.200000 ;
        RECT 6.900000 9.900001 7.300000 10.200000 ;
        RECT 6.900000 8.200000 7.400000 9.900001 ;
        RECT 8.600000 7.900000 9.000000 10.200000 ;
        RECT 12.600000 7.900000 13.000000 10.200000 ;
        RECT 14.200000 8.900001 14.600000 10.200000 ;
        RECT 16.300001 8.000000 16.700001 10.200000 ;
        RECT 22.200001 7.900000 22.600000 10.200000 ;
        RECT 24.600000 7.900000 25.000000 10.200000 ;
        RECT 26.200001 8.900001 26.600000 10.200000 ;
        RECT 27.800001 7.900000 28.200001 10.200000 ;
        RECT 29.400000 8.900001 29.800001 10.200000 ;
        RECT 31.000000 7.900000 31.400000 10.200000 ;
        RECT 33.400002 8.900001 33.799999 10.200000 ;
        RECT 35.000000 7.900000 35.400002 10.200000 ;
        RECT 38.200001 8.900001 38.600002 10.200000 ;
        RECT 39.000000 8.900001 39.400002 10.200000 ;
        RECT 40.600002 8.900001 41.000000 10.200000 ;
        RECT 41.400002 7.900000 41.799999 10.200000 ;
        RECT 44.600002 8.900001 45.000000 10.200000 ;
        RECT 48.600002 8.200000 49.100002 10.200000 ;
        RECT 51.700001 9.900001 52.100002 10.200000 ;
        RECT 51.700001 8.200000 52.200001 9.900001 ;
        RECT 54.200001 8.900001 54.600002 10.200000 ;
        RECT 55.000000 8.900001 55.400002 10.200000 ;
        RECT 56.600002 8.900001 57.000000 10.200000 ;
        RECT 58.299999 9.900001 58.700001 10.200000 ;
        RECT 58.200001 8.200000 58.700001 9.900001 ;
        RECT 61.299999 8.200000 61.799999 10.200000 ;
      LAYER via1 ;
        RECT 46.000000 30.300001 46.400002 30.700001 ;
        RECT 46.500000 30.300001 46.900002 30.700001 ;
        RECT 47.000000 30.300001 47.400002 30.700001 ;
        RECT 47.500000 30.300001 47.900002 30.700001 ;
        RECT 48.000000 30.300001 48.400002 30.700001 ;
        RECT 46.000000 10.300000 46.400002 10.700000 ;
        RECT 46.500000 10.300000 46.900002 10.700000 ;
        RECT 47.000000 10.300000 47.400002 10.700000 ;
        RECT 47.500000 10.300000 47.900002 10.700000 ;
        RECT 48.000000 10.300000 48.400002 10.700000 ;
      LAYER metal2 ;
        RECT 46.900002 30.700001 47.500000 30.800001 ;
        RECT 46.000000 30.300001 48.400002 30.700001 ;
        RECT 46.900002 30.200001 47.500000 30.300001 ;
        RECT 46.900002 10.700000 47.500000 10.800000 ;
        RECT 46.000000 10.300000 48.400002 10.700000 ;
        RECT 46.900002 10.200000 47.500000 10.300000 ;
      LAYER via2 ;
        RECT 46.500000 30.300001 46.900002 30.700001 ;
        RECT 47.000000 30.300001 47.400002 30.700001 ;
        RECT 47.500000 30.300001 47.900002 30.700001 ;
        RECT 48.000000 30.300001 48.400002 30.700001 ;
        RECT 46.500000 10.300000 46.900002 10.700000 ;
        RECT 47.000000 10.300000 47.400002 10.700000 ;
        RECT 47.500000 10.300000 47.900002 10.700000 ;
        RECT 48.000000 10.300000 48.400002 10.700000 ;
      LAYER metal3 ;
        RECT 46.900002 30.700001 47.500000 30.800001 ;
        RECT 46.000000 30.300001 48.400002 30.700001 ;
        RECT 46.900002 30.200001 47.500000 30.300001 ;
        RECT 46.900002 10.700000 47.500000 10.800000 ;
        RECT 46.000000 10.300000 48.400002 10.700000 ;
        RECT 46.900002 10.200000 47.500000 10.300000 ;
      LAYER via3 ;
        RECT 46.100002 30.300001 46.500000 30.700001 ;
        RECT 46.700001 30.300001 47.100002 30.700001 ;
        RECT 47.299999 30.300001 47.700001 30.700001 ;
        RECT 47.900002 30.300001 48.299999 30.700001 ;
        RECT 46.100002 10.300000 46.500000 10.700000 ;
        RECT 46.700001 10.300000 47.100002 10.700000 ;
        RECT 47.299999 10.300000 47.700001 10.700000 ;
        RECT 47.900002 10.300000 48.299999 10.700000 ;
      LAYER metal4 ;
        RECT 46.900002 30.700001 47.500000 30.800001 ;
        RECT 46.000000 30.300001 48.400002 30.700001 ;
        RECT 46.900002 30.200001 47.500000 30.300001 ;
        RECT 46.900002 10.700000 47.500000 10.800000 ;
        RECT 46.000000 10.300000 48.400002 10.700000 ;
        RECT 46.900002 10.200000 47.500000 10.300000 ;
      LAYER via4 ;
        RECT 46.000000 30.300001 46.400002 30.700001 ;
        RECT 46.500000 30.300001 46.900002 30.700001 ;
        RECT 47.000000 30.300001 47.400002 30.700001 ;
        RECT 47.500000 30.300001 47.900002 30.700001 ;
        RECT 48.000000 30.300001 48.400002 30.700001 ;
        RECT 46.000000 10.300000 46.400002 10.700000 ;
        RECT 46.500000 10.300000 46.900002 10.700000 ;
        RECT 47.000000 10.300000 47.400002 10.700000 ;
        RECT 47.500000 10.300000 47.900002 10.700000 ;
        RECT 48.000000 10.300000 48.400002 10.700000 ;
      LAYER metal5 ;
        RECT 46.900002 30.700001 47.500000 30.800001 ;
        RECT 46.000000 30.300001 48.400002 30.700001 ;
        RECT 46.600002 30.200001 47.799999 30.300001 ;
        RECT 46.900002 10.700000 47.500000 10.800000 ;
        RECT 46.000000 10.300000 48.400002 10.700000 ;
        RECT 46.600002 10.200000 47.799999 10.300000 ;
      LAYER via5 ;
        RECT 47.299999 30.200001 47.799999 30.700001 ;
        RECT 47.299999 10.200000 47.799999 10.700000 ;
      LAYER metal6 ;
        RECT 46.000000 -0.600000 48.400002 30.700001 ;
    END
  END gnd
  PIN vdd
    USE POWER ;
    PORT
      LAYER metal1 ;
        RECT 1.400000 20.800001 1.800000 24.500000 ;
        RECT 3.800000 21.100000 4.300000 24.400000 ;
        RECT 3.900000 20.800001 4.300000 21.100000 ;
        RECT 6.900000 20.800001 7.400000 24.400000 ;
        RECT 9.400001 21.100000 9.900001 24.400000 ;
        RECT 9.500000 20.800001 9.900001 21.100000 ;
        RECT 12.500000 20.800001 13.000000 24.400000 ;
        RECT 14.200000 20.800001 14.600000 23.100000 ;
        RECT 15.800000 20.800001 16.200001 23.100000 ;
        RECT 20.600000 20.800001 21.000000 24.500000 ;
        RECT 23.000000 21.100000 23.500000 24.400000 ;
        RECT 23.100000 20.800001 23.500000 21.100000 ;
        RECT 26.100000 20.800001 26.600000 24.400000 ;
        RECT 27.800001 20.800001 28.200001 23.100000 ;
        RECT 29.400000 20.800001 29.800001 25.100000 ;
        RECT 31.800001 20.800001 32.200001 23.100000 ;
        RECT 33.400002 20.800001 33.799999 23.100000 ;
        RECT 35.000000 20.800001 35.400002 23.100000 ;
        RECT 37.400002 20.800001 37.799999 25.100000 ;
        RECT 38.200001 20.800001 38.600002 23.100000 ;
        RECT 39.799999 20.800001 40.200001 23.100000 ;
        RECT 41.400002 20.800001 41.799999 23.100000 ;
        RECT 43.000000 20.800001 43.400002 23.100000 ;
        RECT 44.600002 20.800001 45.100002 24.400000 ;
        RECT 47.700001 21.100000 48.200001 24.400000 ;
        RECT 47.700001 20.800001 48.100002 21.100000 ;
        RECT 52.600002 20.800001 53.100002 24.400000 ;
        RECT 55.700001 21.100000 56.200001 24.400000 ;
        RECT 55.700001 20.800001 56.100002 21.100000 ;
        RECT 58.200001 20.800001 58.600002 23.100000 ;
        RECT 59.799999 20.800001 60.200001 24.500000 ;
        RECT 62.200001 20.800001 62.600002 24.500000 ;
        RECT 0.200000 20.200001 64.599998 20.800001 ;
        RECT 1.400000 16.600000 1.900000 20.200001 ;
        RECT 4.500000 19.900000 4.900000 20.200001 ;
        RECT 4.500000 16.600000 5.000000 19.900000 ;
        RECT 6.200000 17.900000 6.600000 20.200001 ;
        RECT 7.800000 17.900000 8.200000 20.200001 ;
        RECT 11.000000 15.900001 11.400001 20.200001 ;
        RECT 11.800000 17.900000 12.200000 20.200001 ;
        RECT 13.400001 17.900000 13.800000 20.200001 ;
        RECT 14.200000 17.900000 14.600000 20.200001 ;
        RECT 15.800000 17.900000 16.200001 20.200001 ;
        RECT 20.600000 15.900001 21.000000 20.200001 ;
        RECT 21.400000 17.900000 21.800001 20.200001 ;
        RECT 23.000000 17.900000 23.400000 20.200001 ;
        RECT 23.800001 17.900000 24.200001 20.200001 ;
        RECT 25.400000 17.900000 25.800001 20.200001 ;
        RECT 27.000000 17.900000 27.400000 20.200001 ;
        RECT 28.600000 16.600000 29.100000 20.200001 ;
        RECT 31.700001 19.900000 32.100002 20.200001 ;
        RECT 31.700001 16.600000 32.200001 19.900000 ;
        RECT 33.400002 17.900000 33.799999 20.200001 ;
        RECT 35.000000 17.900000 35.400002 20.200001 ;
        RECT 35.799999 17.900000 36.200001 20.200001 ;
        RECT 37.400002 17.900000 37.799999 20.200001 ;
        RECT 39.000000 17.900000 39.400002 20.200001 ;
        RECT 39.799999 17.900000 40.200001 20.200001 ;
        RECT 41.400002 16.100000 41.799999 20.200001 ;
        RECT 43.000000 17.900000 43.400002 20.200001 ;
        RECT 44.600002 17.900000 45.000000 20.200001 ;
        RECT 45.400002 17.900000 45.799999 20.200001 ;
        RECT 47.000000 17.900000 47.400002 20.200001 ;
        RECT 50.200001 17.900000 50.600002 20.200001 ;
        RECT 51.799999 17.900000 52.200001 20.200001 ;
        RECT 53.400002 17.900000 53.799999 20.200001 ;
        RECT 54.200001 17.900000 54.600002 20.200001 ;
        RECT 55.799999 17.900000 56.200001 20.200001 ;
        RECT 57.400002 16.600000 57.900002 20.200001 ;
        RECT 60.500000 19.900000 60.900002 20.200001 ;
        RECT 60.500000 16.600000 61.000000 19.900000 ;
        RECT 63.000000 16.500000 63.400002 20.200001 ;
        RECT 1.400000 0.800000 1.800000 4.500000 ;
        RECT 3.800000 0.800000 4.300000 4.400000 ;
        RECT 6.900000 1.100000 7.400000 4.400000 ;
        RECT 6.900000 0.800000 7.300000 1.100000 ;
        RECT 8.600000 0.800000 9.000000 3.100000 ;
        RECT 10.200000 0.800000 10.600000 3.100000 ;
        RECT 11.000000 0.800000 11.400001 3.100000 ;
        RECT 12.600000 0.800000 13.000000 3.100000 ;
        RECT 14.200000 0.800000 14.600000 3.100000 ;
        RECT 15.000000 0.800000 15.400001 3.100000 ;
        RECT 16.600000 0.800000 17.000000 4.900000 ;
        RECT 20.600000 0.800000 21.000000 3.100000 ;
        RECT 22.200001 0.800000 22.600000 3.100000 ;
        RECT 23.000000 0.800000 23.400000 3.100000 ;
        RECT 24.600000 0.800000 25.000000 3.100000 ;
        RECT 26.200001 0.800000 26.600000 3.100000 ;
        RECT 27.800001 0.800000 28.200001 4.500000 ;
        RECT 29.400000 0.800000 29.800001 3.100000 ;
        RECT 31.000000 0.800000 31.400000 3.100000 ;
        RECT 32.600002 0.800000 33.000000 3.100000 ;
        RECT 33.400002 0.800000 33.799999 3.100000 ;
        RECT 35.000000 0.800000 35.400002 3.100000 ;
        RECT 36.600002 0.800000 37.000000 3.100000 ;
        RECT 38.200001 0.800000 38.600002 3.100000 ;
        RECT 39.000000 0.800000 39.400002 5.100000 ;
        RECT 41.400002 0.800000 41.799999 3.100000 ;
        RECT 43.000000 0.800000 43.400002 3.100000 ;
        RECT 44.600002 0.800000 45.000000 3.100000 ;
        RECT 48.600002 0.800000 49.100002 4.400000 ;
        RECT 51.700001 1.100000 52.200001 4.400000 ;
        RECT 51.700001 0.800000 52.100002 1.100000 ;
        RECT 54.200001 0.800000 54.600002 3.100000 ;
        RECT 55.000000 0.800000 55.400002 5.100000 ;
        RECT 58.200001 1.100000 58.700001 4.400000 ;
        RECT 58.299999 0.800000 58.700001 1.100000 ;
        RECT 61.299999 0.800000 61.799999 4.400000 ;
        RECT 0.200000 0.200000 64.599998 0.800000 ;
      LAYER via1 ;
        RECT 16.400000 20.300001 16.800001 20.700001 ;
        RECT 16.900000 20.300001 17.300001 20.700001 ;
        RECT 17.400000 20.300001 17.800001 20.700001 ;
        RECT 17.900000 20.300001 18.300001 20.700001 ;
        RECT 18.400000 20.300001 18.800001 20.700001 ;
        RECT 16.400000 0.300000 16.800001 0.700000 ;
        RECT 16.900000 0.300000 17.300001 0.700000 ;
        RECT 17.400000 0.300000 17.800001 0.700000 ;
        RECT 17.900000 0.300000 18.300001 0.700000 ;
        RECT 18.400000 0.300000 18.800001 0.700000 ;
      LAYER metal2 ;
        RECT 17.300001 20.700001 17.900000 20.800001 ;
        RECT 16.400000 20.300001 18.800001 20.700001 ;
        RECT 17.300001 20.200001 17.900000 20.300001 ;
        RECT 17.300001 0.700000 17.900000 0.800000 ;
        RECT 16.400000 0.300000 18.800001 0.700000 ;
        RECT 17.300001 0.200000 17.900000 0.300000 ;
      LAYER via2 ;
        RECT 16.900000 20.300001 17.300001 20.700001 ;
        RECT 17.400000 20.300001 17.800001 20.700001 ;
        RECT 17.900000 20.300001 18.300001 20.700001 ;
        RECT 18.400000 20.300001 18.800001 20.700001 ;
        RECT 16.900000 0.300000 17.300001 0.700000 ;
        RECT 17.400000 0.300000 17.800001 0.700000 ;
        RECT 17.900000 0.300000 18.300001 0.700000 ;
        RECT 18.400000 0.300000 18.800001 0.700000 ;
      LAYER metal3 ;
        RECT 17.300001 20.700001 17.900000 20.800001 ;
        RECT 16.400000 20.300001 18.800001 20.700001 ;
        RECT 17.300001 20.200001 17.900000 20.300001 ;
        RECT 17.300001 0.700000 17.900000 0.800000 ;
        RECT 16.400000 0.300000 18.800001 0.700000 ;
        RECT 17.300001 0.200000 17.900000 0.300000 ;
      LAYER via3 ;
        RECT 16.500000 20.300001 16.900000 20.700001 ;
        RECT 17.100000 20.300001 17.500000 20.700001 ;
        RECT 17.700001 20.300001 18.100000 20.700001 ;
        RECT 18.300001 20.300001 18.700001 20.700001 ;
        RECT 16.500000 0.300000 16.900000 0.700000 ;
        RECT 17.100000 0.300000 17.500000 0.700000 ;
        RECT 17.700001 0.300000 18.100000 0.700000 ;
        RECT 18.300001 0.300000 18.700001 0.700000 ;
      LAYER metal4 ;
        RECT 17.300001 20.700001 17.900000 20.800001 ;
        RECT 16.400000 20.300001 18.800001 20.700001 ;
        RECT 17.300001 20.200001 17.900000 20.300001 ;
        RECT 17.300001 0.700000 17.900000 0.800000 ;
        RECT 16.400000 0.300000 18.800001 0.700000 ;
        RECT 17.300001 0.200000 17.900000 0.300000 ;
      LAYER via4 ;
        RECT 16.400000 20.300001 16.800001 20.700001 ;
        RECT 16.900000 20.300001 17.300001 20.700001 ;
        RECT 17.400000 20.300001 17.800001 20.700001 ;
        RECT 17.900000 20.300001 18.300001 20.700001 ;
        RECT 18.400000 20.300001 18.800001 20.700001 ;
        RECT 16.400000 0.300000 16.800001 0.700000 ;
        RECT 16.900000 0.300000 17.300001 0.700000 ;
        RECT 17.400000 0.300000 17.800001 0.700000 ;
        RECT 17.900000 0.300000 18.300001 0.700000 ;
        RECT 18.400000 0.300000 18.800001 0.700000 ;
      LAYER metal5 ;
        RECT 17.300001 20.700001 17.900000 20.800001 ;
        RECT 16.400000 20.300001 18.800001 20.700001 ;
        RECT 17.000000 20.200001 18.200001 20.300001 ;
        RECT 17.300001 0.700000 17.900000 0.800000 ;
        RECT 16.400000 0.300000 18.800001 0.700000 ;
        RECT 17.000000 0.200000 18.200001 0.300000 ;
      LAYER via5 ;
        RECT 17.700001 20.200001 18.200001 20.700001 ;
        RECT 17.700001 0.200000 18.200001 0.700000 ;
      LAYER metal6 ;
        RECT 16.400000 -0.600000 18.800001 30.700001 ;
    END
  END vdd
  PIN s[6]
    PORT
      LAYER metal1 ;
        RECT 19.800001 26.200001 20.200001 29.900000 ;
        RECT 19.800001 25.100000 20.100000 26.200001 ;
        RECT 19.800001 21.100000 20.200001 25.100000 ;
      LAYER via1 ;
        RECT 19.800001 28.800001 20.200001 29.200001 ;
      LAYER metal2 ;
        RECT 21.400000 33.799999 21.800001 34.200001 ;
        RECT 21.400000 30.200001 21.700001 33.799999 ;
        RECT 19.800001 29.800001 20.200001 30.200001 ;
        RECT 21.400000 29.800001 21.800001 30.200001 ;
        RECT 19.800001 29.200001 20.100000 29.800001 ;
        RECT 19.800001 28.800001 20.200001 29.200001 ;
      LAYER metal3 ;
        RECT 19.800001 30.100000 20.200001 30.200001 ;
        RECT 21.400000 30.100000 21.800001 30.200001 ;
        RECT 19.800001 29.800001 21.800001 30.100000 ;
    END
  END s[6]
  PIN s[5]
    PORT
      LAYER metal1 ;
        RECT 0.600000 6.200000 1.000000 9.900001 ;
        RECT 0.600000 5.100000 0.900000 6.200000 ;
        RECT 0.600000 1.100000 1.000000 5.100000 ;
      LAYER via1 ;
        RECT 0.600000 3.800000 1.000000 4.200000 ;
      LAYER metal2 ;
        RECT 0.600000 4.800000 1.000000 5.200000 ;
        RECT 0.600000 4.200000 0.900000 4.800000 ;
        RECT 0.600000 3.800000 1.000000 4.200000 ;
      LAYER metal3 ;
        RECT -2.600000 5.100000 -2.200000 5.200000 ;
        RECT 0.600000 5.100000 1.000000 5.200000 ;
        RECT -2.600000 4.800000 1.000000 5.100000 ;
    END
  END s[5]
  PIN s[4]
    PORT
      LAYER metal1 ;
        RECT 0.600000 26.200001 1.000000 29.900000 ;
        RECT 0.600000 25.100000 0.900000 26.200001 ;
        RECT 0.600000 21.100000 1.000000 25.100000 ;
      LAYER via1 ;
        RECT 0.600000 23.800001 1.000000 24.200001 ;
      LAYER metal2 ;
        RECT 0.600000 24.800001 1.000000 25.200001 ;
        RECT 0.600000 24.200001 0.900000 24.800001 ;
        RECT 0.600000 23.800001 1.000000 24.200001 ;
      LAYER metal3 ;
        RECT -2.600000 25.100000 -2.200000 25.200001 ;
        RECT 0.600000 25.100000 1.000000 25.200001 ;
        RECT -2.600000 24.800001 1.000000 25.100000 ;
    END
  END s[4]
  PIN s[3]
    PORT
      LAYER metal1 ;
        RECT 27.000000 6.200000 27.400000 9.900001 ;
        RECT 27.000000 5.100000 27.300001 6.200000 ;
        RECT 27.000000 1.100000 27.400000 5.100000 ;
      LAYER via1 ;
        RECT 27.000000 1.800000 27.400000 2.200000 ;
      LAYER metal2 ;
        RECT 27.000000 1.800000 27.400000 2.200000 ;
        RECT 27.000000 -1.900000 27.300001 1.800000 ;
        RECT 27.800001 -1.900000 28.200001 -1.800000 ;
        RECT 27.000000 -2.200000 28.200001 -1.900000 ;
    END
  END s[3]
  PIN s[2]
    PORT
      LAYER metal1 ;
        RECT 60.600002 26.200001 61.000000 29.900000 ;
        RECT 60.700001 25.100000 61.000000 26.200001 ;
        RECT 60.600002 21.100000 61.000000 25.100000 ;
      LAYER via1 ;
        RECT 60.600002 28.800001 61.000000 29.200001 ;
      LAYER metal2 ;
        RECT 59.799999 34.100002 60.200001 34.200001 ;
        RECT 59.799999 33.799999 60.900002 34.100002 ;
        RECT 60.600002 29.200001 60.900002 33.799999 ;
        RECT 60.600002 28.800001 61.000000 29.200001 ;
    END
  END s[2]
  PIN s[1]
    PORT
      LAYER metal1 ;
        RECT 63.799999 15.900001 64.200005 19.900000 ;
        RECT 63.900002 14.800000 64.200005 15.900001 ;
        RECT 63.799999 14.100000 64.200005 14.800000 ;
        RECT 64.599998 14.100000 65.000000 14.200000 ;
        RECT 63.799999 13.800000 65.000000 14.100000 ;
        RECT 63.799999 11.100000 64.200005 13.800000 ;
      LAYER via1 ;
        RECT 64.599998 13.800000 65.000000 14.200000 ;
      LAYER metal2 ;
        RECT 64.599998 14.800000 65.000000 15.200000 ;
        RECT 64.599998 14.200000 64.900002 14.800000 ;
        RECT 64.599998 13.800000 65.000000 14.200000 ;
      LAYER metal3 ;
        RECT 64.599998 15.100000 65.000000 15.200000 ;
        RECT 67.000000 15.100000 67.400002 15.200000 ;
        RECT 64.599998 14.800000 67.400002 15.100000 ;
    END
  END s[1]
  PIN s[0]
    PORT
      LAYER metal1 ;
        RECT 63.000000 26.200001 63.400002 29.900000 ;
        RECT 63.100002 25.100000 63.400002 26.200001 ;
        RECT 63.000000 24.100000 63.400002 25.100000 ;
        RECT 64.599998 24.100000 65.000000 24.200001 ;
        RECT 63.000000 23.800001 65.000000 24.100000 ;
        RECT 63.000000 21.100000 63.400002 23.800001 ;
      LAYER via1 ;
        RECT 64.599998 23.800001 65.000000 24.200001 ;
      LAYER metal2 ;
        RECT 64.599998 24.800001 65.000000 25.200001 ;
        RECT 64.599998 24.200001 64.900002 24.800001 ;
        RECT 64.599998 23.800001 65.000000 24.200001 ;
      LAYER metal3 ;
        RECT 64.599998 25.100000 65.000000 25.200001 ;
        RECT 67.000000 25.100000 67.400002 25.200001 ;
        RECT 64.599998 24.800001 67.400002 25.100000 ;
    END
  END s[0]
  PIN x[5]
    PORT
      LAYER metal1 ;
        RECT 0.600000 13.800000 1.400000 14.200000 ;
        RECT 6.200000 12.400001 6.600000 13.200000 ;
      LAYER via1 ;
        RECT 6.200000 12.800000 6.600000 13.200000 ;
      LAYER metal2 ;
        RECT 0.600000 13.800000 1.000000 14.200000 ;
        RECT 0.600000 13.200000 0.900000 13.800000 ;
        RECT 0.600000 12.800000 1.000000 13.200000 ;
        RECT 6.200000 13.100000 6.600000 13.200000 ;
        RECT 7.000000 13.100000 7.400000 13.200000 ;
        RECT 6.200000 12.800000 7.400000 13.100000 ;
      LAYER via2 ;
        RECT 7.000000 12.800000 7.400000 13.200000 ;
      LAYER metal3 ;
        RECT -2.600000 14.100000 -2.200000 14.200000 ;
        RECT 0.600000 14.100000 1.000000 14.200000 ;
        RECT -2.600000 13.800000 1.000000 14.100000 ;
        RECT 0.600000 13.100000 1.000000 13.200000 ;
        RECT 7.000000 13.100000 7.400000 13.200000 ;
        RECT 0.600000 12.800000 7.400000 13.100000 ;
    END
  END x[5]
  PIN x[4]
    PORT
      LAYER metal1 ;
        RECT 14.200000 27.800001 14.600000 28.600000 ;
        RECT 13.000000 27.100000 13.800000 27.200001 ;
        RECT 14.200000 27.100000 14.500000 27.800001 ;
        RECT 13.000000 26.800001 14.500000 27.100000 ;
      LAYER metal2 ;
        RECT 14.200000 33.799999 14.600000 34.200001 ;
        RECT 14.200000 28.200001 14.500000 33.799999 ;
        RECT 14.200000 27.800001 14.600000 28.200001 ;
    END
  END x[4]
  PIN x[3]
    PORT
      LAYER metal1 ;
        RECT 31.800001 27.800001 32.200001 28.600000 ;
        RECT 26.600000 26.800001 27.400000 27.200001 ;
      LAYER via1 ;
        RECT 27.000000 26.800001 27.400000 27.200001 ;
      LAYER metal2 ;
        RECT 31.800001 33.799999 32.200001 34.200001 ;
        RECT 31.800001 28.200001 32.100002 33.799999 ;
        RECT 27.000000 27.800001 27.400000 28.200001 ;
        RECT 31.800001 27.800001 32.200001 28.200001 ;
        RECT 27.000000 27.200001 27.300001 27.800001 ;
        RECT 27.000000 26.800001 27.400000 27.200001 ;
      LAYER metal3 ;
        RECT 27.000000 28.100000 27.400000 28.200001 ;
        RECT 31.800001 28.100000 32.200001 28.200001 ;
        RECT 27.000000 27.800001 32.200001 28.100000 ;
    END
  END x[3]
  PIN x[2]
    PORT
      LAYER metal1 ;
        RECT 43.000000 27.800001 43.400002 28.600000 ;
        RECT 43.000000 27.100000 43.299999 27.800001 ;
        RECT 43.799999 27.100000 44.600002 27.200001 ;
        RECT 43.000000 26.800001 44.600002 27.100000 ;
      LAYER via1 ;
        RECT 43.799999 26.800001 44.200001 27.200001 ;
      LAYER metal2 ;
        RECT 43.799999 33.799999 44.200001 34.200001 ;
        RECT 43.799999 27.200001 44.100002 33.799999 ;
        RECT 43.799999 26.800001 44.200001 27.200001 ;
    END
  END x[2]
  PIN x[1]
    PORT
      LAYER metal1 ;
        RECT 44.600002 8.100000 45.000000 8.600000 ;
        RECT 44.600002 7.800000 47.299999 8.100000 ;
        RECT 47.000000 7.100000 47.299999 7.800000 ;
        RECT 47.799999 7.100000 48.600002 7.200000 ;
        RECT 47.000000 6.800000 48.600002 7.100000 ;
        RECT 47.799999 6.100000 48.100002 6.800000 ;
        RECT 49.400002 6.100000 49.799999 6.200000 ;
        RECT 47.799999 5.800000 49.799999 6.100000 ;
      LAYER via1 ;
        RECT 49.400002 5.800000 49.799999 6.200000 ;
      LAYER metal2 ;
        RECT 49.400002 5.800000 49.799999 6.200000 ;
        RECT 49.400002 -1.800000 49.700001 5.800000 ;
        RECT 49.400002 -2.200000 49.799999 -1.800000 ;
    END
  END x[1]
  PIN x[0]
    PORT
      LAYER metal1 ;
        RECT 58.200001 27.800001 58.600002 28.600000 ;
        RECT 61.799999 7.100000 62.600002 7.200000 ;
        RECT 63.000000 7.100000 63.400002 7.200000 ;
        RECT 61.799999 6.800000 63.400002 7.100000 ;
      LAYER via1 ;
        RECT 63.000000 6.800000 63.400002 7.200000 ;
      LAYER metal2 ;
        RECT 58.200001 27.800001 58.600002 28.200001 ;
        RECT 58.200001 27.100000 58.500000 27.800001 ;
        RECT 58.200001 26.800001 59.299999 27.100000 ;
        RECT 59.000000 18.200001 59.299999 26.800001 ;
        RECT 59.000000 17.800001 59.400002 18.200001 ;
        RECT 63.000000 17.800001 63.400002 18.200001 ;
        RECT 63.000000 7.200000 63.299999 17.800001 ;
        RECT 63.000000 6.800000 63.400002 7.200000 ;
      LAYER metal3 ;
        RECT 59.000000 18.100000 59.400002 18.200001 ;
        RECT 63.000000 18.100000 63.400002 18.200001 ;
        RECT 67.000000 18.100000 67.400002 18.200001 ;
        RECT 59.000000 17.800001 67.400002 18.100000 ;
    END
  END x[0]
  PIN y[5]
    PORT
      LAYER metal1 ;
        RECT 3.600000 14.300000 4.000000 14.400001 ;
        RECT 3.600000 14.200000 5.000000 14.300000 ;
        RECT 3.600000 14.000000 5.800000 14.200000 ;
        RECT 4.700000 13.900001 5.800000 14.000000 ;
        RECT 5.000000 13.800000 5.800000 13.900001 ;
        RECT 7.800000 12.400001 8.200000 13.200000 ;
      LAYER via1 ;
        RECT 5.400000 13.800000 5.800000 14.200000 ;
        RECT 7.800000 12.800000 8.200000 13.200000 ;
      LAYER metal2 ;
        RECT 5.400000 15.800000 5.800000 16.200001 ;
        RECT 5.400000 14.200000 5.700000 15.800000 ;
        RECT 5.400000 14.100000 5.800000 14.200000 ;
        RECT 6.200000 14.100000 6.600000 14.200000 ;
        RECT 5.400000 13.800000 6.600000 14.100000 ;
        RECT 7.800000 13.800000 8.200000 14.200000 ;
        RECT 7.800000 13.200000 8.100000 13.800000 ;
        RECT 7.800000 12.800000 8.200000 13.200000 ;
      LAYER via2 ;
        RECT 6.200000 13.800000 6.600000 14.200000 ;
      LAYER metal3 ;
        RECT -2.600000 16.100000 -2.200000 16.200001 ;
        RECT 5.400000 16.100000 5.800000 16.200001 ;
        RECT -2.600000 15.800000 5.800000 16.100000 ;
        RECT 6.200000 14.100000 6.600000 14.200000 ;
        RECT 7.800000 14.100000 8.200000 14.200000 ;
        RECT 6.200000 13.800000 8.200000 14.100000 ;
    END
  END y[5]
  PIN y[4]
    PORT
      LAYER metal1 ;
        RECT 15.800000 27.800001 16.200001 28.600000 ;
        RECT 8.600000 27.100000 9.400001 27.200001 ;
        RECT 8.600000 27.000000 9.700000 27.100000 ;
        RECT 8.600000 26.800001 10.800000 27.000000 ;
        RECT 9.400001 26.700001 10.800000 26.800001 ;
        RECT 10.400001 26.600000 10.800000 26.700001 ;
      LAYER metal2 ;
        RECT 19.800001 33.799999 20.200001 34.200001 ;
        RECT 19.800001 31.200001 20.100000 33.799999 ;
        RECT 8.600000 30.800001 9.000000 31.200001 ;
        RECT 15.800000 30.800001 16.200001 31.200001 ;
        RECT 19.800001 30.800001 20.200001 31.200001 ;
        RECT 8.600000 27.200001 8.900001 30.800001 ;
        RECT 15.800000 28.200001 16.100000 30.800001 ;
        RECT 15.800000 27.800001 16.200001 28.200001 ;
        RECT 8.600000 26.800001 9.000000 27.200001 ;
      LAYER metal3 ;
        RECT 8.600000 31.100000 9.000000 31.200001 ;
        RECT 15.800000 31.100000 16.200001 31.200001 ;
        RECT 19.800001 31.100000 20.200001 31.200001 ;
        RECT 8.600000 30.800001 20.200001 31.100000 ;
    END
  END y[4]
  PIN y[3]
    PORT
      LAYER metal1 ;
        RECT 27.800001 27.800001 28.200001 28.600000 ;
        RECT 22.200001 27.100000 23.000000 27.200001 ;
        RECT 22.200001 27.000000 23.300001 27.100000 ;
        RECT 22.200001 26.800001 24.400000 27.000000 ;
        RECT 23.000000 26.700001 24.400000 26.800001 ;
        RECT 24.000000 26.600000 24.400000 26.700001 ;
      LAYER metal2 ;
        RECT 27.800001 33.799999 28.200001 34.200001 ;
        RECT 27.800001 28.200001 28.100000 33.799999 ;
        RECT 22.200001 27.800001 22.600000 28.200001 ;
        RECT 27.800001 27.800001 28.200001 28.200001 ;
        RECT 22.200001 27.200001 22.500000 27.800001 ;
        RECT 27.800001 27.200001 28.100000 27.800001 ;
        RECT 22.200001 26.800001 22.600000 27.200001 ;
        RECT 27.800001 26.800001 28.200001 27.200001 ;
      LAYER metal3 ;
        RECT 22.200001 27.800001 22.600000 28.200001 ;
        RECT 22.200001 27.100000 22.500000 27.800001 ;
        RECT 27.800001 27.100000 28.200001 27.200001 ;
        RECT 22.200001 26.800001 28.200001 27.100000 ;
    END
  END y[3]
  PIN y[2]
    PORT
      LAYER metal1 ;
        RECT 41.400002 27.800001 41.799999 28.600000 ;
        RECT 48.200001 27.100000 49.000000 27.200001 ;
        RECT 47.900002 27.000000 49.000000 27.100000 ;
        RECT 46.799999 26.800001 49.000000 27.000000 ;
        RECT 46.799999 26.700001 48.200001 26.800001 ;
        RECT 46.799999 26.600000 47.200001 26.700001 ;
      LAYER via1 ;
        RECT 48.600002 26.800001 49.000000 27.200001 ;
      LAYER metal2 ;
        RECT 41.400002 33.799999 41.799999 34.200001 ;
        RECT 41.400002 28.200001 41.700001 33.799999 ;
        RECT 41.400002 27.800001 41.799999 28.200001 ;
        RECT 48.600002 27.800001 49.000000 28.200001 ;
        RECT 41.400002 27.200001 41.700001 27.800001 ;
        RECT 48.600002 27.200001 48.900002 27.800001 ;
        RECT 41.400002 26.800001 41.799999 27.200001 ;
        RECT 48.600002 26.800001 49.000000 27.200001 ;
      LAYER metal3 ;
        RECT 48.600002 27.800001 49.000000 28.200001 ;
        RECT 41.400002 27.100000 41.799999 27.200001 ;
        RECT 48.600002 27.100000 48.900002 27.800001 ;
        RECT 41.400002 26.800001 48.900002 27.100000 ;
    END
  END y[2]
  PIN y[1]
    PORT
      LAYER metal1 ;
        RECT 38.200001 7.800000 38.600002 8.600000 ;
        RECT 52.200001 7.100000 53.000000 7.200000 ;
        RECT 51.900002 7.000000 53.000000 7.100000 ;
        RECT 50.799999 6.800000 53.000000 7.000000 ;
        RECT 50.799999 6.700000 52.200001 6.800000 ;
        RECT 50.799999 6.600000 51.200001 6.700000 ;
      LAYER via1 ;
        RECT 52.600002 6.800000 53.000000 7.200000 ;
      LAYER metal2 ;
        RECT 38.200001 8.100000 38.600002 8.200000 ;
        RECT 39.000000 8.100000 39.400002 8.200000 ;
        RECT 38.200001 7.800000 39.400002 8.100000 ;
        RECT 52.600002 7.800000 53.000000 8.200000 ;
        RECT 52.600002 7.200000 52.900002 7.800000 ;
        RECT 52.600002 6.800000 53.000000 7.200000 ;
        RECT 52.600002 1.200000 52.900002 6.800000 ;
        RECT 51.000000 0.800000 51.400002 1.200000 ;
        RECT 52.600002 0.800000 53.000000 1.200000 ;
        RECT 51.000000 -1.800000 51.299999 0.800000 ;
        RECT 51.000000 -2.200000 51.400002 -1.800000 ;
      LAYER via2 ;
        RECT 39.000000 7.800000 39.400002 8.200000 ;
      LAYER metal3 ;
        RECT 39.000000 8.100000 39.400002 8.200000 ;
        RECT 52.600002 8.100000 53.000000 8.200000 ;
        RECT 38.200001 7.800000 53.000000 8.100000 ;
        RECT 51.000000 1.100000 51.400002 1.200000 ;
        RECT 52.600002 1.100000 53.000000 1.200000 ;
        RECT 51.000000 0.800000 53.000000 1.100000 ;
    END
  END y[1]
  PIN y[0]
    PORT
      LAYER metal1 ;
        RECT 54.200001 7.800000 54.600002 8.600000 ;
        RECT 57.400002 7.100000 58.200001 7.200000 ;
        RECT 57.400002 7.000000 58.500000 7.100000 ;
        RECT 57.400002 6.800000 59.600002 7.000000 ;
        RECT 58.200001 6.700000 59.600002 6.800000 ;
        RECT 59.200001 6.600000 59.600002 6.700000 ;
      LAYER metal2 ;
        RECT 54.200001 7.800000 54.600002 8.200000 ;
        RECT 54.200001 7.200000 54.500000 7.800000 ;
        RECT 54.200001 6.800000 54.600002 7.200000 ;
        RECT 56.600002 7.100000 57.000000 7.200000 ;
        RECT 57.400002 7.100000 57.799999 7.200000 ;
        RECT 56.600002 6.800000 57.799999 7.100000 ;
        RECT 57.400002 1.200000 57.700001 6.800000 ;
        RECT 57.400002 0.800000 57.799999 1.200000 ;
        RECT 59.000000 0.800000 59.400002 1.200000 ;
        RECT 59.000000 -1.800000 59.299999 0.800000 ;
        RECT 59.000000 -2.200000 59.400002 -1.800000 ;
      LAYER metal3 ;
        RECT 54.200001 7.100000 54.600002 7.200000 ;
        RECT 56.600002 7.100000 57.000000 7.200000 ;
        RECT 54.200001 6.800000 57.000000 7.100000 ;
        RECT 57.400002 1.100000 57.799999 1.200000 ;
        RECT 59.000000 1.100000 59.400002 1.200000 ;
        RECT 57.400002 0.800000 59.400002 1.100000 ;
    END
  END y[0]
  OBS
      LAYER metal1 ;
        RECT 2.200000 27.600000 2.600000 29.900000 ;
        RECT 3.000000 27.900000 3.400000 29.900000 ;
        RECT 5.200000 28.100000 6.000000 29.900000 ;
        RECT 3.000000 27.600000 4.300000 27.900000 ;
        RECT 1.500000 27.300001 2.600000 27.600000 ;
        RECT 3.900000 27.500000 4.300000 27.600000 ;
        RECT 4.600000 27.400000 5.400000 27.800001 ;
        RECT 1.500000 25.800001 1.800000 27.300001 ;
        RECT 3.000000 27.100000 3.800000 27.200001 ;
        RECT 5.700000 27.100000 6.000000 28.100000 ;
        RECT 7.800000 27.900000 8.200000 29.900000 ;
        RECT 6.300000 27.400000 6.700000 27.800001 ;
        RECT 7.000000 27.600000 8.200000 27.900000 ;
        RECT 8.600000 27.900000 9.000000 29.900000 ;
        RECT 10.800000 29.200001 11.600000 29.900000 ;
        RECT 10.200000 28.800001 11.600000 29.200001 ;
        RECT 10.800000 28.100000 11.600000 28.800001 ;
        RECT 8.600000 27.600000 9.900001 27.900000 ;
        RECT 7.000000 27.500000 7.400000 27.600000 ;
        RECT 9.500000 27.500000 9.900001 27.600000 ;
        RECT 10.200000 27.400000 11.000000 27.800001 ;
        RECT 3.000000 27.000000 4.100000 27.100000 ;
        RECT 3.000000 26.800001 5.200000 27.000000 ;
        RECT 3.800000 26.700001 5.200000 26.800001 ;
        RECT 4.800000 26.600000 5.200000 26.700001 ;
        RECT 5.500000 26.800001 6.000000 27.100000 ;
        RECT 6.400000 27.200001 6.700000 27.400000 ;
        RECT 6.400000 26.800001 6.800000 27.200001 ;
        RECT 7.400000 26.800001 8.200000 27.200001 ;
        RECT 11.300000 27.100000 11.600000 28.100000 ;
        RECT 13.400001 27.900000 13.800000 29.900000 ;
        RECT 11.900001 27.400000 12.300000 27.800001 ;
        RECT 12.600000 27.600000 13.800000 27.900000 ;
        RECT 12.600000 27.500000 13.000000 27.600000 ;
        RECT 11.100000 26.800001 11.600000 27.100000 ;
        RECT 12.000000 27.200001 12.300000 27.400000 ;
        RECT 12.000000 26.800001 12.400001 27.200001 ;
        RECT 2.200000 25.800001 2.600000 26.600000 ;
        RECT 5.500000 26.200001 5.800000 26.800001 ;
        RECT 11.100000 26.200001 11.400001 26.800001 ;
        RECT 4.100000 26.100000 4.500000 26.200001 ;
        RECT 4.100000 25.800001 4.900000 26.100000 ;
        RECT 5.400000 25.800001 5.800000 26.200001 ;
        RECT 9.700000 26.100000 10.100000 26.200001 ;
        RECT 9.700000 25.800001 10.500000 26.100000 ;
        RECT 11.000000 25.800001 11.400001 26.200001 ;
        RECT 1.200000 25.400000 1.800000 25.800001 ;
        RECT 4.500000 25.700001 4.900000 25.800001 ;
        RECT 1.500000 25.100000 1.800000 25.400000 ;
        RECT 5.500000 25.100000 5.800000 25.800001 ;
        RECT 10.100000 25.700001 10.500000 25.800001 ;
        RECT 11.100000 25.100000 11.400001 25.800001 ;
        RECT 1.500000 24.800001 2.600000 25.100000 ;
        RECT 2.200000 21.100000 2.600000 24.800001 ;
        RECT 3.000000 24.800001 4.300000 25.100000 ;
        RECT 3.000000 21.100000 3.400000 24.800001 ;
        RECT 3.900000 24.700001 4.300000 24.800001 ;
        RECT 5.200000 21.100000 6.000000 25.100000 ;
        RECT 7.000000 24.800001 8.200000 25.100000 ;
        RECT 7.000000 24.700001 7.400000 24.800001 ;
        RECT 7.800000 21.100000 8.200000 24.800001 ;
        RECT 8.600000 24.800001 9.900001 25.100000 ;
        RECT 8.600000 21.100000 9.000000 24.800001 ;
        RECT 9.500000 24.700001 9.900001 24.800001 ;
        RECT 10.800000 21.100000 11.600000 25.100000 ;
        RECT 12.600000 24.800001 13.800000 25.100000 ;
        RECT 12.600000 24.700001 13.000000 24.800001 ;
        RECT 13.400001 21.100000 13.800000 24.800001 ;
        RECT 14.200000 24.100000 14.600000 24.200001 ;
        RECT 15.000000 24.100000 15.400001 29.900000 ;
        RECT 14.200000 23.800001 15.400001 24.100000 ;
        RECT 15.000000 21.100000 15.400001 23.800001 ;
        RECT 16.600000 22.100000 17.000000 29.900000 ;
        RECT 21.400000 27.600000 21.800001 29.900000 ;
        RECT 22.200001 27.900000 22.600000 29.900000 ;
        RECT 24.400000 28.100000 25.200001 29.900000 ;
        RECT 22.200001 27.600000 23.500000 27.900000 ;
        RECT 20.700001 27.300001 21.800001 27.600000 ;
        RECT 23.100000 27.500000 23.500000 27.600000 ;
        RECT 23.800001 27.400000 24.600000 27.800001 ;
        RECT 20.700001 25.800001 21.000000 27.300001 ;
        RECT 24.900000 27.100000 25.200001 28.100000 ;
        RECT 27.000000 27.900000 27.400000 29.900000 ;
        RECT 25.500000 27.400000 25.900000 27.800001 ;
        RECT 26.200001 27.600000 27.400000 27.900000 ;
        RECT 28.600000 28.100000 29.000000 29.900000 ;
        RECT 30.200001 28.900000 30.600000 29.900000 ;
        RECT 29.400000 28.100000 29.800001 28.600000 ;
        RECT 28.600000 27.800001 29.800001 28.100000 ;
        RECT 26.200001 27.500000 26.600000 27.600000 ;
        RECT 24.700001 26.800001 25.200001 27.100000 ;
        RECT 25.600000 27.200001 25.900000 27.400000 ;
        RECT 25.600000 26.800001 26.000000 27.200001 ;
        RECT 28.600000 27.100000 29.000000 27.800001 ;
        RECT 30.300001 27.200001 30.600000 28.900000 ;
        RECT 28.600000 26.800001 29.700001 27.100000 ;
        RECT 30.200001 26.800001 30.600000 27.200001 ;
        RECT 21.400000 25.800001 21.800001 26.600000 ;
        RECT 24.700001 26.200001 25.000000 26.800001 ;
        RECT 23.300001 26.100000 23.700001 26.200001 ;
        RECT 23.300001 25.800001 24.100000 26.100000 ;
        RECT 24.600000 25.800001 25.000000 26.200001 ;
        RECT 20.400000 25.400000 21.000000 25.800001 ;
        RECT 23.700001 25.700001 24.100000 25.800001 ;
        RECT 20.700001 25.100000 21.000000 25.400000 ;
        RECT 24.700001 25.100000 25.000000 25.800001 ;
        RECT 20.700001 24.800001 21.800001 25.100000 ;
        RECT 18.200001 22.100000 18.600000 22.200001 ;
        RECT 16.600000 21.800001 18.600000 22.100000 ;
        RECT 16.600000 21.100000 17.000000 21.800001 ;
        RECT 21.400000 21.100000 21.800001 24.800001 ;
        RECT 22.200001 24.800001 23.500000 25.100000 ;
        RECT 22.200001 21.100000 22.600000 24.800001 ;
        RECT 23.100000 24.700001 23.500000 24.800001 ;
        RECT 24.400000 22.200001 25.200001 25.100000 ;
        RECT 26.200001 24.800001 27.400000 25.100000 ;
        RECT 26.200001 24.700001 26.600000 24.800001 ;
        RECT 24.400000 21.800001 25.800001 22.200001 ;
        RECT 24.400000 21.100000 25.200001 21.800001 ;
        RECT 27.000000 21.100000 27.400000 24.800001 ;
        RECT 28.600000 21.100000 29.000000 26.800001 ;
        RECT 29.400000 26.200001 29.700001 26.800001 ;
        RECT 29.400000 25.800001 29.800001 26.200001 ;
        RECT 30.300001 25.100000 30.600000 26.800001 ;
        RECT 31.000000 26.100000 31.400000 26.200001 ;
        RECT 32.600002 26.100000 33.000000 29.900000 ;
        RECT 33.700001 28.200001 34.100002 29.900000 ;
        RECT 36.600002 28.900000 37.000000 29.900000 ;
        RECT 33.700001 27.900000 34.600002 28.200001 ;
        RECT 31.000000 25.800001 33.000000 26.100000 ;
        RECT 33.400002 26.100000 33.799999 26.200001 ;
        RECT 34.200001 26.100000 34.600002 27.900000 ;
        RECT 35.000000 26.800001 35.400002 27.600000 ;
        RECT 36.600002 27.200001 36.900002 28.900000 ;
        RECT 37.400002 27.800001 37.799999 28.600000 ;
        RECT 38.500000 28.200001 38.900002 29.900000 ;
        RECT 38.500000 27.900000 39.400002 28.200001 ;
        RECT 36.600002 26.800001 37.000000 27.200001 ;
        RECT 33.400002 25.800001 34.600002 26.100000 ;
        RECT 31.000000 25.400000 31.400000 25.800001 ;
        RECT 32.600002 25.100000 33.000000 25.800001 ;
        RECT 33.400002 25.100000 33.799999 25.200001 ;
        RECT 30.200001 24.700001 31.100000 25.100000 ;
        RECT 30.700001 22.200001 31.100000 24.700001 ;
        RECT 30.200001 21.800001 31.100000 22.200001 ;
        RECT 30.700001 21.100000 31.100000 21.800001 ;
        RECT 32.600002 24.800001 33.799999 25.100000 ;
        RECT 32.600002 21.100000 33.000000 24.800001 ;
        RECT 33.400002 24.400000 33.799999 24.800001 ;
        RECT 34.200001 21.100000 34.600002 25.800001 ;
        RECT 35.799999 25.400000 36.200001 26.200001 ;
        RECT 36.600002 25.100000 36.900002 26.800001 ;
        RECT 36.100002 24.700001 37.000000 25.100000 ;
        RECT 36.100002 22.200001 36.500000 24.700001 ;
        RECT 38.200001 24.400000 38.600002 25.200001 ;
        RECT 35.799999 21.800001 36.500000 22.200001 ;
        RECT 36.100002 21.100000 36.500000 21.800001 ;
        RECT 39.000000 24.100000 39.400002 27.900000 ;
        RECT 39.799999 27.100000 40.200001 27.600000 ;
        RECT 40.600002 27.100000 41.000000 29.900000 ;
        RECT 39.799999 26.800001 41.000000 27.100000 ;
        RECT 39.799999 24.100000 40.200001 24.200001 ;
        RECT 39.000000 23.800001 40.200001 24.100000 ;
        RECT 39.000000 21.100000 39.400002 23.800001 ;
        RECT 40.600002 21.100000 41.000000 26.800001 ;
        RECT 41.400002 25.800001 41.799999 26.200001 ;
        RECT 41.400002 25.100000 41.700001 25.800001 ;
        RECT 42.200001 25.100000 42.600002 29.900000 ;
        RECT 43.799999 27.900000 44.200001 29.900000 ;
        RECT 46.000000 28.100000 46.799999 29.900000 ;
        RECT 43.799999 27.600000 45.000000 27.900000 ;
        RECT 44.600002 27.500000 45.000000 27.600000 ;
        RECT 45.299999 27.400000 45.700001 27.800001 ;
        RECT 45.299999 27.200001 45.600002 27.400000 ;
        RECT 45.200001 26.800001 45.600002 27.200001 ;
        RECT 46.000000 27.100000 46.299999 28.100000 ;
        RECT 48.600002 27.900000 49.000000 29.900000 ;
        RECT 46.600002 27.400000 47.400002 27.800001 ;
        RECT 47.700001 27.600000 49.000000 27.900000 ;
        RECT 51.799999 27.900000 52.200001 29.900000 ;
        RECT 54.000000 28.100000 54.799999 29.900000 ;
        RECT 51.799999 27.600000 53.000000 27.900000 ;
        RECT 47.700001 27.500000 48.100002 27.600000 ;
        RECT 52.600002 27.500000 53.000000 27.600000 ;
        RECT 53.299999 27.400000 53.700001 27.800001 ;
        RECT 53.299999 27.200001 53.600002 27.400000 ;
        RECT 46.000000 26.800001 46.500000 27.100000 ;
        RECT 51.799999 26.800001 52.600002 27.200001 ;
        RECT 53.200001 26.800001 53.600002 27.200001 ;
        RECT 54.000000 27.100000 54.299999 28.100000 ;
        RECT 56.600002 27.900000 57.000000 29.900000 ;
        RECT 54.600002 27.400000 55.400002 27.800001 ;
        RECT 55.700001 27.600000 57.000000 27.900000 ;
        RECT 55.700001 27.500000 56.100002 27.600000 ;
        RECT 56.200001 27.100000 57.000000 27.200001 ;
        RECT 54.000000 26.800001 54.500000 27.100000 ;
        RECT 55.900002 27.000000 57.000000 27.100000 ;
        RECT 46.200001 26.200001 46.500000 26.800001 ;
        RECT 54.200001 26.200001 54.500000 26.800001 ;
        RECT 54.799999 26.800001 57.000000 27.000000 ;
        RECT 54.799999 26.700001 56.200001 26.800001 ;
        RECT 54.799999 26.600000 55.200001 26.700001 ;
        RECT 45.400002 26.100000 45.799999 26.200001 ;
        RECT 46.200001 26.100000 46.600002 26.200001 ;
        RECT 47.500000 26.100000 47.900002 26.200001 ;
        RECT 45.400002 25.800001 46.600002 26.100000 ;
        RECT 47.100002 25.800001 47.900002 26.100000 ;
        RECT 54.200001 25.800001 54.600002 26.200001 ;
        RECT 55.500000 26.100000 55.900002 26.200001 ;
        RECT 55.100002 25.800001 55.900002 26.100000 ;
        RECT 46.200001 25.100000 46.500000 25.800001 ;
        RECT 47.100002 25.700001 47.500000 25.800001 ;
        RECT 54.200001 25.100000 54.500000 25.800001 ;
        RECT 55.100002 25.700001 55.500000 25.800001 ;
        RECT 41.400002 24.800001 42.600002 25.100000 ;
        RECT 42.200001 21.100000 42.600002 24.800001 ;
        RECT 43.799999 24.800001 45.000000 25.100000 ;
        RECT 43.799999 21.100000 44.200001 24.800001 ;
        RECT 44.600002 24.700001 45.000000 24.800001 ;
        RECT 46.000000 21.100000 46.799999 25.100000 ;
        RECT 47.700001 24.800001 49.000000 25.100000 ;
        RECT 47.700001 24.700001 48.100002 24.800001 ;
        RECT 48.600002 21.100000 49.000000 24.800001 ;
        RECT 51.799999 24.800001 53.000000 25.100000 ;
        RECT 51.799999 21.100000 52.200001 24.800001 ;
        RECT 52.600002 24.700001 53.000000 24.800001 ;
        RECT 54.000000 21.100000 54.799999 25.100000 ;
        RECT 55.700001 24.800001 57.000000 25.100000 ;
        RECT 55.700001 24.700001 56.100002 24.800001 ;
        RECT 56.600002 21.100000 57.000000 24.800001 ;
        RECT 57.400002 21.100000 57.799999 29.900000 ;
        RECT 59.000000 27.600000 59.400002 29.900000 ;
        RECT 61.400002 27.600000 61.799999 29.900000 ;
        RECT 59.000000 27.300001 60.100002 27.600000 ;
        RECT 61.400002 27.300001 62.500000 27.600000 ;
        RECT 59.000000 26.100000 59.400002 26.600000 ;
        RECT 58.200001 25.800001 59.400002 26.100000 ;
        RECT 59.799999 25.800001 60.100002 27.300001 ;
        RECT 61.400002 25.800001 61.799999 26.600000 ;
        RECT 62.200001 25.800001 62.500000 27.300001 ;
        RECT 58.200001 25.200001 58.500000 25.800001 ;
        RECT 59.799999 25.400000 60.400002 25.800001 ;
        RECT 62.200001 25.400000 62.799999 25.800001 ;
        RECT 58.200001 24.800001 58.600002 25.200001 ;
        RECT 59.799999 25.100000 60.100002 25.400000 ;
        RECT 62.200001 25.100000 62.500000 25.400000 ;
        RECT 59.000000 24.800001 60.100002 25.100000 ;
        RECT 61.400002 24.800001 62.500000 25.100000 ;
        RECT 59.000000 21.100000 59.400002 24.800001 ;
        RECT 61.400002 21.100000 61.799999 24.800001 ;
        RECT 0.600000 16.200001 1.000000 19.900000 ;
        RECT 1.400000 16.200001 1.800000 16.300001 ;
        RECT 0.600000 15.900001 1.800000 16.200001 ;
        RECT 2.800000 15.900001 3.600000 19.900000 ;
        RECT 4.500000 16.200001 4.900000 16.300001 ;
        RECT 5.400000 16.200001 5.800000 19.900000 ;
        RECT 4.500000 15.900001 5.800000 16.200001 ;
        RECT 3.000000 15.200000 3.300000 15.900001 ;
        RECT 3.900000 15.200000 4.300000 15.300000 ;
        RECT 3.000000 14.800000 3.400000 15.200000 ;
        RECT 3.900000 14.900001 4.700000 15.200000 ;
        RECT 4.300000 14.800000 4.700000 14.900001 ;
        RECT 7.000000 15.100000 7.400000 19.900000 ;
        RECT 7.800000 15.800000 8.200000 16.200001 ;
        RECT 7.800000 15.100000 8.100000 15.800000 ;
        RECT 7.000000 14.800000 8.100000 15.100000 ;
        RECT 3.000000 14.200000 3.300000 14.800000 ;
        RECT 2.000000 13.800000 2.400000 14.200000 ;
        RECT 2.100000 13.600000 2.400000 13.800000 ;
        RECT 2.800000 13.900001 3.300000 14.200000 ;
        RECT 1.400000 13.400001 1.800000 13.500000 ;
        RECT 0.600000 13.100000 1.800000 13.400001 ;
        RECT 2.100000 13.200000 2.500000 13.600000 ;
        RECT 0.600000 11.100000 1.000000 13.100000 ;
        RECT 2.800000 12.900001 3.100000 13.900001 ;
        RECT 3.400000 13.200000 4.200000 13.600000 ;
        RECT 4.500000 13.400001 4.900000 13.500000 ;
        RECT 4.500000 13.100000 5.800000 13.400001 ;
        RECT 2.800000 11.100000 3.600000 12.900001 ;
        RECT 5.400000 11.100000 5.800000 13.100000 ;
        RECT 7.000000 11.100000 7.400000 14.800000 ;
        RECT 8.600000 13.100000 9.000000 19.900000 ;
        RECT 9.700000 16.300001 10.100000 19.900000 ;
        RECT 9.700000 15.900001 10.600000 16.300001 ;
        RECT 9.400001 14.800000 9.800000 15.600000 ;
        RECT 10.200000 14.200000 10.500000 15.900001 ;
        RECT 9.400001 13.800000 9.800000 14.200000 ;
        RECT 10.200000 13.800000 10.600000 14.200000 ;
        RECT 11.800000 14.100000 12.200000 14.200000 ;
        RECT 11.000000 13.800000 12.200000 14.100000 ;
        RECT 9.400001 13.100000 9.700000 13.800000 ;
        RECT 8.600000 12.800000 9.700000 13.100000 ;
        RECT 8.600000 11.100000 9.000000 12.800000 ;
        RECT 10.200000 12.200000 10.500000 13.800000 ;
        RECT 11.000000 13.200000 11.300000 13.800000 ;
        RECT 11.800000 13.400001 12.200000 13.800000 ;
        RECT 11.000000 12.400001 11.400001 13.200000 ;
        RECT 12.600000 13.100000 13.000000 19.900000 ;
        RECT 13.400001 15.800000 13.800000 16.600000 ;
        RECT 14.200000 15.800000 14.600000 16.600000 ;
        RECT 15.000000 13.100000 15.400001 19.900000 ;
        RECT 19.300001 16.300001 19.700001 19.900000 ;
        RECT 19.300001 15.900001 20.200001 16.300001 ;
        RECT 19.000000 14.800000 19.400000 15.600000 ;
        RECT 19.800001 14.200000 20.100000 15.900001 ;
        RECT 15.800000 13.400001 16.200001 14.200000 ;
        RECT 19.800001 14.100000 20.200001 14.200000 ;
        RECT 21.400000 14.100000 21.800001 14.200000 ;
        RECT 19.800001 13.800000 21.800001 14.100000 ;
        RECT 12.600000 12.800000 13.500000 13.100000 ;
        RECT 13.100000 12.200000 13.500000 12.800000 ;
        RECT 14.500000 12.800000 15.400001 13.100000 ;
        RECT 14.500000 12.200000 14.900001 12.800000 ;
        RECT 19.800001 12.200000 20.100000 13.800000 ;
        RECT 21.400000 13.400001 21.800001 13.800000 ;
        RECT 20.600000 12.400001 21.000000 13.200000 ;
        RECT 22.200001 13.100000 22.600000 19.900000 ;
        RECT 23.000000 15.800000 23.400000 16.600000 ;
        RECT 24.600000 14.100000 25.000000 19.900000 ;
        RECT 25.400000 14.100000 25.800001 14.200000 ;
        RECT 24.600000 13.800000 25.800001 14.100000 ;
        RECT 22.200001 12.800000 23.100000 13.100000 ;
        RECT 10.200000 11.100000 10.600000 12.200000 ;
        RECT 13.100000 11.800000 13.800000 12.200000 ;
        RECT 14.500000 11.800000 15.400001 12.200000 ;
        RECT 13.100000 11.100000 13.500000 11.800000 ;
        RECT 14.500000 11.100000 14.900001 11.800000 ;
        RECT 19.800001 11.100000 20.200001 12.200000 ;
        RECT 22.700001 11.100000 23.100000 12.800000 ;
        RECT 23.800001 12.400001 24.200001 13.200000 ;
        RECT 24.600000 11.100000 25.000000 13.800000 ;
        RECT 25.400000 13.400001 25.800001 13.800000 ;
        RECT 26.200001 13.100000 26.600000 19.900000 ;
        RECT 27.000000 15.800000 27.400000 16.600000 ;
        RECT 27.800001 16.200001 28.200001 19.900000 ;
        RECT 28.600000 16.200001 29.000000 16.300001 ;
        RECT 27.800001 15.900001 29.000000 16.200001 ;
        RECT 30.000000 15.900001 30.800001 19.900000 ;
        RECT 31.700001 16.200001 32.100002 16.300001 ;
        RECT 32.600002 16.200001 33.000000 19.900000 ;
        RECT 31.700001 15.900001 33.000000 16.200001 ;
        RECT 30.200001 15.200000 30.500000 15.900001 ;
        RECT 33.400002 15.800000 33.799999 16.600000 ;
        RECT 31.100000 15.200000 31.500000 15.300000 ;
        RECT 30.200001 14.800000 30.600000 15.200000 ;
        RECT 31.100000 14.900001 31.900000 15.200000 ;
        RECT 31.500000 14.800000 31.900000 14.900001 ;
        RECT 30.200001 14.200000 30.500000 14.800000 ;
        RECT 27.800001 13.800000 28.600000 14.200000 ;
        RECT 29.200001 13.800000 29.600000 14.200000 ;
        RECT 29.300001 13.600000 29.600000 13.800000 ;
        RECT 30.000000 13.900001 30.500000 14.200000 ;
        RECT 30.800001 14.300000 31.200001 14.400001 ;
        RECT 30.800001 14.200000 32.200001 14.300000 ;
        RECT 30.800001 14.000000 33.000000 14.200000 ;
        RECT 31.900000 13.900001 33.000000 14.000000 ;
        RECT 28.600000 13.400001 29.000000 13.500000 ;
        RECT 27.800001 13.100000 29.000000 13.400001 ;
        RECT 29.300001 13.200000 29.700001 13.600000 ;
        RECT 26.200001 12.800000 27.100000 13.100000 ;
        RECT 26.700001 12.200000 27.100000 12.800000 ;
        RECT 26.200001 11.800000 27.100000 12.200000 ;
        RECT 26.700001 11.100000 27.100000 11.800000 ;
        RECT 27.800001 11.100000 28.200001 13.100000 ;
        RECT 30.000000 12.900001 30.300001 13.900001 ;
        RECT 32.200001 13.800000 33.000000 13.900001 ;
        RECT 30.600000 13.200000 31.400000 13.600000 ;
        RECT 31.700001 13.400001 32.100002 13.500000 ;
        RECT 31.700001 13.100000 33.000000 13.400001 ;
        RECT 34.200001 13.100000 34.600002 19.900000 ;
        RECT 35.000000 14.100000 35.400002 14.200000 ;
        RECT 35.799999 14.100000 36.200001 14.200000 ;
        RECT 35.000000 13.800000 36.200001 14.100000 ;
        RECT 36.600002 14.100000 37.000000 19.900000 ;
        RECT 37.400002 14.100000 37.799999 14.200000 ;
        RECT 36.600002 13.800000 37.799999 14.100000 ;
        RECT 35.000000 13.400001 35.400002 13.800000 ;
        RECT 30.000000 11.100000 30.800001 12.900001 ;
        RECT 32.600002 11.100000 33.000000 13.100000 ;
        RECT 33.700001 12.800000 34.600002 13.100000 ;
        RECT 33.700001 12.200000 34.100002 12.800000 ;
        RECT 35.799999 12.400001 36.200001 13.200000 ;
        RECT 33.400002 11.800000 34.100002 12.200000 ;
        RECT 33.700001 11.100000 34.100002 11.800000 ;
        RECT 36.600002 11.100000 37.000000 13.800000 ;
        RECT 37.400002 13.400001 37.799999 13.800000 ;
        RECT 38.200001 13.100000 38.600002 19.900000 ;
        RECT 40.600002 17.900000 41.000000 19.900000 ;
        RECT 39.000000 15.800000 39.400002 16.600000 ;
        RECT 40.700001 15.800000 41.000000 17.900000 ;
        RECT 42.200001 15.900001 42.600002 19.900000 ;
        RECT 40.700001 15.500000 41.900002 15.800000 ;
        RECT 40.600002 14.800000 41.000000 15.200000 ;
        RECT 39.799999 13.800000 40.200001 14.600000 ;
        RECT 40.700001 14.400001 41.000000 14.800000 ;
        RECT 40.700001 14.100000 41.200001 14.400001 ;
        RECT 40.799999 14.000000 41.200001 14.100000 ;
        RECT 41.600002 13.800000 41.900002 15.500000 ;
        RECT 42.299999 15.200000 42.600002 15.900001 ;
        RECT 43.000000 15.800000 43.400002 16.600000 ;
        RECT 42.200001 14.800000 42.600002 15.200000 ;
        RECT 43.799999 15.100000 44.200001 19.900000 ;
        RECT 45.400002 15.800000 45.799999 16.600000 ;
        RECT 41.600002 13.700000 42.000000 13.800000 ;
        RECT 40.500000 13.500000 42.000000 13.700000 ;
        RECT 39.900002 13.400001 42.000000 13.500000 ;
        RECT 39.900002 13.200000 40.799999 13.400001 ;
        RECT 39.900002 13.100000 40.200001 13.200000 ;
        RECT 42.299999 13.100000 42.600002 14.800000 ;
        RECT 43.000000 14.800000 44.200001 15.100000 ;
        RECT 43.000000 14.200000 43.299999 14.800000 ;
        RECT 43.000000 13.800000 43.400002 14.200000 ;
        RECT 43.799999 13.100000 44.200001 14.800000 ;
        RECT 44.600002 13.400001 45.000000 14.200000 ;
        RECT 46.200001 13.100000 46.600002 19.900000 ;
        RECT 47.000000 13.400001 47.400002 14.200000 ;
        RECT 51.000000 14.100000 51.400002 19.900000 ;
        RECT 51.799999 14.100000 52.200001 14.200000 ;
        RECT 51.000000 13.800000 52.200001 14.100000 ;
        RECT 38.200001 12.800000 39.100002 13.100000 ;
        RECT 38.700001 11.100000 39.100002 12.800000 ;
        RECT 39.799999 11.100000 40.200001 13.100000 ;
        RECT 41.900002 12.600000 42.600002 13.100000 ;
        RECT 43.299999 12.800000 44.200001 13.100000 ;
        RECT 45.700001 12.800000 46.600002 13.100000 ;
        RECT 41.900002 11.100000 42.299999 12.600000 ;
        RECT 43.299999 11.100000 43.700001 12.800000 ;
        RECT 45.700001 12.200000 46.100002 12.800000 ;
        RECT 50.200001 12.400001 50.600002 13.200000 ;
        RECT 45.400002 11.800000 46.100002 12.200000 ;
        RECT 45.700001 11.100000 46.100002 11.800000 ;
        RECT 51.000000 11.100000 51.400002 13.800000 ;
        RECT 51.799999 13.400001 52.200001 13.800000 ;
        RECT 52.600002 14.100000 53.000000 19.900000 ;
        RECT 53.400002 15.800000 53.799999 16.600000 ;
        RECT 54.200001 15.800000 54.600002 16.600000 ;
        RECT 53.400002 15.100000 53.700001 15.800000 ;
        RECT 55.000000 15.100000 55.400002 19.900000 ;
        RECT 56.600002 16.200001 57.000000 19.900000 ;
        RECT 57.400002 16.200001 57.799999 16.300001 ;
        RECT 56.600002 15.900001 57.799999 16.200001 ;
        RECT 58.799999 15.900001 59.600002 19.900000 ;
        RECT 60.500000 16.200001 60.900002 16.300001 ;
        RECT 61.400002 16.200001 61.799999 19.900000 ;
        RECT 60.500000 15.900001 61.799999 16.200001 ;
        RECT 62.200001 16.200001 62.600002 19.900000 ;
        RECT 62.200001 15.900001 63.299999 16.200001 ;
        RECT 53.400002 14.800000 55.400002 15.100000 ;
        RECT 53.400002 14.100000 53.799999 14.200000 ;
        RECT 52.600002 13.800000 53.799999 14.100000 ;
        RECT 52.600002 13.100000 53.000000 13.800000 ;
        RECT 55.000000 13.100000 55.400002 14.800000 ;
        RECT 59.000000 15.800000 59.400002 15.900001 ;
        RECT 59.000000 15.200000 59.299999 15.800000 ;
        RECT 63.000000 15.600000 63.299999 15.900001 ;
        RECT 59.900002 15.200000 60.299999 15.300000 ;
        RECT 63.000000 15.200000 63.600002 15.600000 ;
        RECT 59.000000 14.800000 59.400002 15.200000 ;
        RECT 59.900002 14.900001 60.700001 15.200000 ;
        RECT 60.299999 14.800000 60.700001 14.900001 ;
        RECT 59.000000 14.200000 59.299999 14.800000 ;
        RECT 62.200001 14.400001 62.600002 15.200000 ;
        RECT 55.799999 13.400001 56.200001 14.200000 ;
        RECT 56.600002 13.800000 57.400002 14.200000 ;
        RECT 58.000000 13.800000 58.400002 14.200000 ;
        RECT 58.100002 13.600000 58.400002 13.800000 ;
        RECT 58.799999 13.900001 59.299999 14.200000 ;
        RECT 59.600002 14.300000 60.000000 14.400001 ;
        RECT 59.600002 14.200000 61.000000 14.300000 ;
        RECT 59.600002 14.000000 61.799999 14.200000 ;
        RECT 60.700001 13.900001 61.799999 14.000000 ;
        RECT 57.400002 13.400001 57.799999 13.500000 ;
        RECT 52.600002 12.800000 53.500000 13.100000 ;
        RECT 53.100002 11.100000 53.500000 12.800000 ;
        RECT 54.500000 12.800000 55.400002 13.100000 ;
        RECT 56.600002 13.100000 57.799999 13.400001 ;
        RECT 58.100002 13.200000 58.500000 13.600000 ;
        RECT 54.500000 11.100000 54.900002 12.800000 ;
        RECT 56.600002 11.100000 57.000000 13.100000 ;
        RECT 58.799999 12.900001 59.100002 13.900001 ;
        RECT 61.000000 13.800000 61.799999 13.900001 ;
        RECT 63.000000 13.700000 63.299999 15.200000 ;
        RECT 59.400002 13.200000 60.200001 13.600000 ;
        RECT 60.500000 13.400001 60.900002 13.500000 ;
        RECT 62.200001 13.400001 63.299999 13.700000 ;
        RECT 60.500000 13.100000 61.799999 13.400001 ;
        RECT 58.799999 11.100000 59.600002 12.900001 ;
        RECT 61.400002 11.100000 61.799999 13.100000 ;
        RECT 62.200001 11.100000 62.600002 13.400001 ;
        RECT 2.200000 7.600000 2.600000 9.900001 ;
        RECT 3.000000 7.900000 3.400000 9.900001 ;
        RECT 5.200000 8.100000 6.000000 9.900001 ;
        RECT 3.000000 7.600000 4.200000 7.900000 ;
        RECT 1.500000 7.300000 2.600000 7.600000 ;
        RECT 3.800000 7.500000 4.200000 7.600000 ;
        RECT 4.500000 7.400000 4.900000 7.800000 ;
        RECT 1.500000 5.800000 1.800000 7.300000 ;
        RECT 4.500000 7.200000 4.800000 7.400000 ;
        RECT 3.000000 6.800000 3.800000 7.200000 ;
        RECT 4.400000 6.800000 4.800000 7.200000 ;
        RECT 5.200000 7.100000 5.500000 8.100000 ;
        RECT 7.800000 7.900000 8.200000 9.900001 ;
        RECT 9.900001 8.200000 10.300000 9.900001 ;
        RECT 5.800000 7.400000 6.600000 7.800000 ;
        RECT 6.900000 7.600000 8.200000 7.900000 ;
        RECT 9.400001 7.900000 10.300000 8.200000 ;
        RECT 11.300000 8.200000 11.700000 9.900001 ;
        RECT 11.300000 7.900000 12.200000 8.200000 ;
        RECT 6.900000 7.500000 7.300000 7.600000 ;
        RECT 7.400000 7.100000 8.200000 7.200000 ;
        RECT 5.200000 6.800000 5.700000 7.100000 ;
        RECT 7.100000 7.000000 8.200000 7.100000 ;
        RECT 2.200000 6.100000 2.600000 6.600000 ;
        RECT 5.400000 6.200000 5.700000 6.800000 ;
        RECT 6.000000 6.800000 8.200000 7.000000 ;
        RECT 8.600000 6.800000 9.000000 7.600000 ;
        RECT 6.000000 6.700000 7.400000 6.800000 ;
        RECT 6.000000 6.600000 6.400000 6.700000 ;
        RECT 5.400000 6.100000 5.800000 6.200000 ;
        RECT 6.700000 6.100000 7.100000 6.200000 ;
        RECT 2.200000 5.800000 5.800000 6.100000 ;
        RECT 6.300000 5.800000 7.100000 6.100000 ;
        RECT 9.400001 6.100000 9.800000 7.900000 ;
        RECT 11.000000 7.100000 11.400001 7.200000 ;
        RECT 11.800000 7.100000 12.200000 7.900000 ;
        RECT 11.000000 6.800000 12.200000 7.100000 ;
        RECT 12.600000 7.100000 13.000000 7.600000 ;
        RECT 13.400001 7.100000 13.800000 9.900001 ;
        RECT 14.200000 7.800000 14.600000 8.600000 ;
        RECT 15.000000 7.900000 15.400001 9.900001 ;
        RECT 17.100000 8.400001 17.500000 9.900001 ;
        RECT 17.100000 7.900000 17.800001 8.400001 ;
        RECT 20.900000 8.200000 21.300001 9.900001 ;
        RECT 23.300001 9.200000 23.700001 9.900001 ;
        RECT 23.000000 8.800000 23.700001 9.200000 ;
        RECT 23.300001 8.200000 23.700001 8.800000 ;
        RECT 20.900000 7.900000 21.800001 8.200000 ;
        RECT 23.300001 7.900000 24.200001 8.200000 ;
        RECT 15.100000 7.800000 15.400001 7.900000 ;
        RECT 15.100000 7.600000 16.000000 7.800000 ;
        RECT 15.100000 7.500000 17.200001 7.600000 ;
        RECT 15.700000 7.300000 17.200001 7.500000 ;
        RECT 16.800001 7.200000 17.200001 7.300000 ;
        RECT 12.600000 6.800000 13.800000 7.100000 ;
        RECT 14.200000 7.100000 14.600000 7.200000 ;
        RECT 15.000000 7.100000 15.400001 7.200000 ;
        RECT 14.200000 6.800000 15.400001 7.100000 ;
        RECT 16.000000 6.900000 16.400000 7.000000 ;
        RECT 9.400001 5.800000 11.300000 6.100000 ;
        RECT 1.200000 5.400000 1.800000 5.800000 ;
        RECT 1.500000 5.100000 1.800000 5.400000 ;
        RECT 5.400000 5.100000 5.700000 5.800000 ;
        RECT 6.300000 5.700000 6.700000 5.800000 ;
        RECT 1.500000 4.800000 2.600000 5.100000 ;
        RECT 2.200000 1.100000 2.600000 4.800000 ;
        RECT 3.000000 4.800000 4.200000 5.100000 ;
        RECT 3.000000 1.100000 3.400000 4.800000 ;
        RECT 3.800000 4.700000 4.200000 4.800000 ;
        RECT 5.200000 1.100000 6.000000 5.100000 ;
        RECT 6.900000 4.800000 8.200000 5.100000 ;
        RECT 6.900000 4.700000 7.300000 4.800000 ;
        RECT 7.800000 1.100000 8.200000 4.800000 ;
        RECT 9.400001 1.100000 9.800000 5.800000 ;
        RECT 11.000000 5.200000 11.300000 5.800000 ;
        RECT 10.200000 4.400000 10.600000 5.200000 ;
        RECT 11.000000 4.400000 11.400001 5.200000 ;
        RECT 11.800000 1.100000 12.200000 6.800000 ;
        RECT 13.400001 1.100000 13.800000 6.800000 ;
        RECT 15.000000 6.400000 15.400001 6.800000 ;
        RECT 15.900001 6.600000 16.400000 6.900000 ;
        RECT 15.900001 6.200000 16.200001 6.600000 ;
        RECT 15.800000 5.800000 16.200001 6.200000 ;
        RECT 16.800001 5.500000 17.100000 7.200000 ;
        RECT 17.500000 6.200000 17.800001 7.900000 ;
        RECT 17.400000 5.800000 17.800001 6.200000 ;
        RECT 15.900001 5.200000 17.100000 5.500000 ;
        RECT 15.900001 3.100000 16.200001 5.200000 ;
        RECT 17.500000 5.100000 17.800001 5.800000 ;
        RECT 20.600000 5.100000 21.000000 5.200000 ;
        RECT 15.800000 1.100000 16.200001 3.100000 ;
        RECT 17.400000 4.800000 21.000000 5.100000 ;
        RECT 17.400000 1.100000 17.800001 4.800000 ;
        RECT 20.600000 4.400000 21.000000 4.800000 ;
        RECT 21.400000 5.100000 21.800001 7.900000 ;
        RECT 22.200001 6.800000 22.600000 7.600000 ;
        RECT 23.000000 5.100000 23.400000 5.200000 ;
        RECT 21.400000 4.800000 23.400000 5.100000 ;
        RECT 21.400000 1.100000 21.800001 4.800000 ;
        RECT 23.000000 4.400000 23.400000 4.800000 ;
        RECT 23.800001 1.100000 24.200001 7.900000 ;
        RECT 24.600000 7.100000 25.000000 7.600000 ;
        RECT 25.400000 7.100000 25.800001 9.900001 ;
        RECT 26.200001 7.800000 26.600000 8.600000 ;
        RECT 28.600000 7.600000 29.000000 9.900001 ;
        RECT 29.400000 7.800000 29.800001 8.600000 ;
        RECT 24.600000 6.800000 25.800001 7.100000 ;
        RECT 25.400000 1.100000 25.800001 6.800000 ;
        RECT 27.900000 7.300000 29.000000 7.600000 ;
        RECT 27.900000 5.800000 28.200001 7.300000 ;
        RECT 30.200001 7.100000 30.600000 9.900001 ;
        RECT 32.299999 8.200000 32.700001 9.900001 ;
        RECT 31.800001 8.100000 32.700001 8.200000 ;
        RECT 33.400002 8.100000 33.799999 8.600000 ;
        RECT 31.800001 7.800000 33.799999 8.100000 ;
        RECT 31.000000 7.100000 31.400000 7.600000 ;
        RECT 30.200001 6.800000 31.400000 7.100000 ;
        RECT 28.600000 6.100000 29.000000 6.600000 ;
        RECT 29.400000 6.100000 29.800001 6.200000 ;
        RECT 28.600000 5.800000 29.800001 6.100000 ;
        RECT 27.600000 5.400000 28.200001 5.800000 ;
        RECT 27.900000 5.100000 28.200001 5.400000 ;
        RECT 27.900000 4.800000 29.000000 5.100000 ;
        RECT 28.600000 1.100000 29.000000 4.800000 ;
        RECT 30.200001 1.100000 30.600000 6.800000 ;
        RECT 31.800001 1.100000 32.200001 7.800000 ;
        RECT 34.200001 7.100000 34.600002 9.900001 ;
        RECT 36.299999 8.200000 36.700001 9.900001 ;
        RECT 35.799999 7.900000 36.700001 8.200000 ;
        RECT 35.000000 7.100000 35.400002 7.600000 ;
        RECT 34.200001 6.800000 35.400002 7.100000 ;
        RECT 32.600002 5.100000 33.000000 5.200000 ;
        RECT 33.400002 5.100000 33.799999 5.200000 ;
        RECT 32.600002 4.800000 33.799999 5.100000 ;
        RECT 32.600002 4.400000 33.000000 4.800000 ;
        RECT 34.200001 1.100000 34.600002 6.800000 ;
        RECT 35.799999 1.100000 36.200001 7.900000 ;
        RECT 37.400002 7.100000 37.799999 9.900001 ;
        RECT 39.799999 8.800000 40.200001 9.900001 ;
        RECT 39.000000 7.800000 39.400002 8.600000 ;
        RECT 39.000000 7.100000 39.299999 7.800000 ;
        RECT 39.900002 7.200000 40.200001 8.800000 ;
        RECT 42.700001 9.200000 43.100002 9.900001 ;
        RECT 42.700001 8.800000 43.400002 9.200000 ;
        RECT 42.700001 8.200000 43.100002 8.800000 ;
        RECT 42.200001 7.900000 43.100002 8.200000 ;
        RECT 37.400002 6.800000 39.299999 7.100000 ;
        RECT 39.799999 6.800000 40.200001 7.200000 ;
        RECT 41.400002 6.800000 41.799999 7.600000 ;
        RECT 36.600002 4.400000 37.000000 5.200000 ;
        RECT 37.400002 1.100000 37.799999 6.800000 ;
        RECT 39.000000 6.200000 39.299999 6.800000 ;
        RECT 39.000000 5.800000 39.400002 6.200000 ;
        RECT 39.900002 5.100000 40.200001 6.800000 ;
        RECT 40.600002 5.400000 41.000000 6.200000 ;
        RECT 39.799999 4.700000 40.700001 5.100000 ;
        RECT 40.299999 1.100000 40.700001 4.700000 ;
        RECT 42.200001 1.100000 42.600002 7.900000 ;
        RECT 43.000000 6.800000 43.400002 7.200000 ;
        RECT 43.000000 6.100000 43.299999 6.800000 ;
        RECT 43.799999 6.100000 44.200001 9.900001 ;
        RECT 47.799999 7.900000 48.200001 9.900001 ;
        RECT 50.000000 9.200000 50.799999 9.900001 ;
        RECT 50.000000 8.800000 51.400002 9.200000 ;
        RECT 50.000000 8.100000 50.799999 8.800000 ;
        RECT 47.799999 7.600000 49.000000 7.900000 ;
        RECT 48.600002 7.500000 49.000000 7.600000 ;
        RECT 49.299999 7.400000 49.700001 7.800000 ;
        RECT 49.299999 7.200000 49.600002 7.400000 ;
        RECT 49.200001 6.800000 49.600002 7.200000 ;
        RECT 50.000000 7.100000 50.299999 8.100000 ;
        RECT 52.600002 7.900000 53.000000 9.900001 ;
        RECT 50.600002 7.400000 51.400002 7.800000 ;
        RECT 51.700001 7.600000 53.000000 7.900000 ;
        RECT 51.700001 7.500000 52.100002 7.600000 ;
        RECT 53.400002 7.100000 53.799999 9.900001 ;
        RECT 55.799999 8.800000 56.200001 9.900001 ;
        RECT 55.000000 7.800000 55.400002 8.600000 ;
        RECT 55.000000 7.100000 55.299999 7.800000 ;
        RECT 55.900002 7.200000 56.200001 8.800000 ;
        RECT 57.400002 7.900000 57.799999 9.900001 ;
        RECT 59.600002 8.100000 60.400002 9.900001 ;
        RECT 57.400002 7.600000 58.700001 7.900000 ;
        RECT 58.299999 7.500000 58.700001 7.600000 ;
        RECT 59.000000 7.400000 59.799999 7.800000 ;
        RECT 50.000000 6.800000 50.500000 7.100000 ;
        RECT 43.000000 5.800000 44.200001 6.100000 ;
        RECT 43.000000 5.100000 43.400002 5.200000 ;
        RECT 43.799999 5.100000 44.200001 5.800000 ;
        RECT 50.200001 6.200000 50.500000 6.800000 ;
        RECT 53.400002 6.800000 55.299999 7.100000 ;
        RECT 55.799999 6.800000 56.200001 7.200000 ;
        RECT 60.100002 7.100000 60.400002 8.100000 ;
        RECT 62.200001 7.900000 62.600002 9.900001 ;
        RECT 60.700001 7.400000 61.100002 7.800000 ;
        RECT 61.400002 7.600000 62.600002 7.900000 ;
        RECT 61.400002 7.500000 61.799999 7.600000 ;
        RECT 50.200001 5.800000 50.600002 6.200000 ;
        RECT 51.500000 6.100000 51.900002 6.200000 ;
        RECT 51.100002 5.800000 51.900002 6.100000 ;
        RECT 50.200001 5.100000 50.500000 5.800000 ;
        RECT 51.100002 5.700000 51.500000 5.800000 ;
        RECT 43.000000 4.800000 44.200001 5.100000 ;
        RECT 43.000000 4.400000 43.400002 4.800000 ;
        RECT 43.799999 1.100000 44.200001 4.800000 ;
        RECT 47.799999 4.800000 49.000000 5.100000 ;
        RECT 47.799999 1.100000 48.200001 4.800000 ;
        RECT 48.600002 4.700000 49.000000 4.800000 ;
        RECT 50.000000 1.100000 50.799999 5.100000 ;
        RECT 51.700001 4.800000 53.000000 5.100000 ;
        RECT 51.700001 4.700000 52.100002 4.800000 ;
        RECT 52.600002 1.100000 53.000000 4.800000 ;
        RECT 53.400002 1.100000 53.799999 6.800000 ;
        RECT 55.900002 5.100000 56.200001 6.800000 ;
        RECT 59.900002 6.800000 60.400002 7.100000 ;
        RECT 60.799999 7.200000 61.100002 7.400000 ;
        RECT 60.799999 6.800000 61.200001 7.200000 ;
        RECT 59.900002 6.200000 60.200001 6.800000 ;
        RECT 56.600002 5.400000 57.000000 6.200000 ;
        RECT 58.500000 6.100000 58.900002 6.200000 ;
        RECT 58.500000 5.800000 59.299999 6.100000 ;
        RECT 59.799999 5.800000 60.200001 6.200000 ;
        RECT 58.900002 5.700000 59.299999 5.800000 ;
        RECT 59.900002 5.100000 60.200001 5.800000 ;
        RECT 55.799999 4.700000 56.700001 5.100000 ;
        RECT 56.299999 1.100000 56.700001 4.700000 ;
        RECT 57.400002 4.800000 58.700001 5.100000 ;
        RECT 57.400002 1.100000 57.799999 4.800000 ;
        RECT 58.299999 4.700000 58.700001 4.800000 ;
        RECT 59.600002 1.100000 60.400002 5.100000 ;
        RECT 61.400002 4.800000 62.600002 5.100000 ;
        RECT 61.400002 4.700000 61.799999 4.800000 ;
        RECT 62.200001 1.100000 62.600002 4.800000 ;
      LAYER via1 ;
        RECT 7.800000 26.800001 8.200000 27.200001 ;
        RECT 18.200001 21.800001 18.600000 22.200001 ;
        RECT 25.400000 21.800001 25.800001 22.200001 ;
        RECT 35.799999 25.800001 36.200001 26.200001 ;
        RECT 38.200001 24.800001 38.600002 25.200001 ;
        RECT 39.799999 23.800001 40.200001 24.200001 ;
        RECT 47.000000 27.400000 47.400002 27.800001 ;
        RECT 55.000000 27.400000 55.400002 27.800001 ;
        RECT 56.600002 26.800001 57.000000 27.200001 ;
        RECT 57.400002 21.800001 57.799999 22.200001 ;
        RECT 1.400000 15.900001 1.800000 16.300001 ;
        RECT 1.400000 13.100000 1.800000 13.500000 ;
        RECT 3.800000 13.200000 4.200000 13.600000 ;
        RECT 3.000000 11.800000 3.400000 12.200000 ;
        RECT 11.000000 12.800000 11.400001 13.200000 ;
        RECT 22.200001 15.800000 22.600000 16.200001 ;
        RECT 15.800000 13.800000 16.200001 14.200000 ;
        RECT 20.600000 12.800000 21.000000 13.200000 ;
        RECT 10.200000 11.800000 10.600000 12.200000 ;
        RECT 13.400001 11.800000 13.800000 12.200000 ;
        RECT 15.000000 11.800000 15.400001 12.200000 ;
        RECT 19.800001 11.800000 20.200001 12.200000 ;
        RECT 23.800001 12.800000 24.200001 13.200000 ;
        RECT 28.600000 15.900001 29.000000 16.300001 ;
        RECT 28.600000 13.100000 29.000000 13.500000 ;
        RECT 32.600002 13.800000 33.000000 14.200000 ;
        RECT 31.000000 13.200000 31.400000 13.600000 ;
        RECT 35.799999 13.800000 36.200001 14.200000 ;
        RECT 30.200001 11.800000 30.600000 12.200000 ;
        RECT 35.799999 12.800000 36.200001 13.200000 ;
        RECT 42.200001 16.800001 42.600002 17.200001 ;
        RECT 44.600002 13.800000 45.000000 14.200000 ;
        RECT 47.000000 13.800000 47.400002 14.200000 ;
        RECT 50.200001 12.800000 50.600002 13.200000 ;
        RECT 57.400002 15.900001 57.799999 16.300001 ;
        RECT 53.400002 13.800000 53.799999 14.200000 ;
        RECT 62.200001 14.800000 62.600002 15.200000 ;
        RECT 55.799999 13.800000 56.200001 14.200000 ;
        RECT 57.400002 13.100000 57.799999 13.500000 ;
        RECT 61.400002 13.800000 61.799999 14.200000 ;
        RECT 59.799999 13.200000 60.200001 13.600000 ;
        RECT 6.200000 7.400000 6.600000 7.800000 ;
        RECT 7.800000 6.800000 8.200000 7.200000 ;
        RECT 10.200000 4.800000 10.600000 5.200000 ;
        RECT 29.400000 5.800000 29.800001 6.200000 ;
        RECT 35.799999 6.800000 36.200001 7.200000 ;
        RECT 33.400002 4.800000 33.799999 5.200000 ;
        RECT 43.000000 8.800000 43.400002 9.200000 ;
        RECT 36.600002 4.800000 37.000000 5.200000 ;
        RECT 40.600002 5.800000 41.000000 6.200000 ;
        RECT 51.000000 8.800000 51.400002 9.200000 ;
        RECT 51.000000 7.400000 51.400002 7.800000 ;
        RECT 59.799999 8.800000 60.200001 9.200000 ;
        RECT 56.600002 5.800000 57.000000 6.200000 ;
      LAYER metal2 ;
        RECT 7.800000 28.800001 8.200000 29.200001 ;
        RECT 10.200000 29.100000 10.600000 29.200001 ;
        RECT 11.000000 29.100000 11.400001 29.200001 ;
        RECT 10.200000 28.800001 11.400001 29.100000 ;
        RECT 3.900000 27.800001 4.300000 27.900000 ;
        RECT 3.900000 27.500000 6.700000 27.800001 ;
        RECT 7.000000 27.500000 7.400000 27.900000 ;
        RECT 3.000000 26.800001 3.400000 27.200001 ;
        RECT 1.400000 26.100000 1.800000 26.200001 ;
        RECT 2.200000 26.100000 2.600000 26.200001 ;
        RECT 1.400000 25.800001 2.600000 26.100000 ;
        RECT 3.000000 25.200001 3.300000 26.800001 ;
        RECT 3.000000 24.800001 3.400000 25.200001 ;
        RECT 3.900000 25.100000 4.200000 27.500000 ;
        RECT 4.600000 27.400000 5.000000 27.500000 ;
        RECT 6.300000 27.400000 6.700000 27.500000 ;
        RECT 7.100000 27.100000 7.400000 27.500000 ;
        RECT 4.600000 26.800001 7.400000 27.100000 ;
        RECT 7.800000 27.200001 8.100000 28.800001 ;
        RECT 37.400002 28.100000 37.799999 28.200001 ;
        RECT 38.200001 28.100000 38.600002 28.200001 ;
        RECT 9.500000 27.800001 9.900001 27.900000 ;
        RECT 9.500000 27.500000 12.300000 27.800001 ;
        RECT 12.600000 27.500000 13.000000 27.900000 ;
        RECT 7.800000 26.800001 8.200000 27.200001 ;
        RECT 4.600000 26.100000 4.900000 26.800001 ;
        RECT 4.500000 25.700001 4.900000 26.100000 ;
        RECT 5.400000 25.800001 5.800000 26.200001 ;
        RECT 5.400000 25.200001 5.700000 25.800001 ;
        RECT 3.900000 24.700001 4.300000 25.100000 ;
        RECT 5.400000 24.800001 5.800000 25.200001 ;
        RECT 7.100000 25.100000 7.400000 26.800001 ;
        RECT 7.000000 24.700001 7.400000 25.100000 ;
        RECT 9.500000 25.100000 9.800000 27.500000 ;
        RECT 10.200000 27.400000 10.600000 27.500000 ;
        RECT 11.900001 27.400000 12.300000 27.500000 ;
        RECT 12.700000 27.100000 13.000000 27.500000 ;
        RECT 10.200000 26.800001 13.000000 27.100000 ;
        RECT 10.200000 26.100000 10.500000 26.800001 ;
        RECT 10.100000 25.700001 10.500000 26.100000 ;
        RECT 12.700000 25.100000 13.000000 26.800001 ;
        RECT 23.100000 27.800001 23.500000 27.900000 ;
        RECT 23.100000 27.500000 25.900000 27.800001 ;
        RECT 26.200001 27.500000 26.600000 27.900000 ;
        RECT 37.400002 27.800001 38.600002 28.100000 ;
        RECT 39.799999 27.800001 40.200001 28.200001 ;
        RECT 9.500000 24.700001 9.900001 25.100000 ;
        RECT 12.600000 24.700001 13.000000 25.100000 ;
        RECT 21.400000 25.800001 21.800001 26.200001 ;
        RECT 14.200000 23.800001 14.600000 24.200001 ;
        RECT 1.400000 15.900001 1.800000 16.300001 ;
        RECT 4.500000 15.900001 4.900000 16.300001 ;
        RECT 14.200000 16.200001 14.500000 23.800001 ;
        RECT 18.200001 22.100000 18.600000 22.200001 ;
        RECT 19.000000 22.100000 19.400000 22.200001 ;
        RECT 18.200001 21.800001 19.400000 22.100000 ;
        RECT 20.600000 21.800001 21.000000 22.200001 ;
        RECT 1.400000 14.200000 1.700000 15.900001 ;
        RECT 3.900000 14.900001 4.300000 15.300000 ;
        RECT 3.900000 14.200000 4.200000 14.900001 ;
        RECT 1.400000 13.900001 4.200000 14.200000 ;
        RECT 1.400000 13.500000 1.700000 13.900001 ;
        RECT 2.100000 13.500000 2.500000 13.600000 ;
        RECT 3.800000 13.500000 4.200000 13.600000 ;
        RECT 4.600000 13.500000 4.900000 15.900001 ;
        RECT 7.800000 15.800000 8.200000 16.200001 ;
        RECT 13.400001 15.800000 13.800000 16.200001 ;
        RECT 14.200000 15.800000 14.600000 16.200001 ;
        RECT 7.800000 15.200000 8.100000 15.800000 ;
        RECT 13.400001 15.200000 13.700000 15.800000 ;
        RECT 14.200000 15.200000 14.500000 15.800000 ;
        RECT 7.800000 14.800000 8.200000 15.200000 ;
        RECT 8.600000 15.100000 9.000000 15.200000 ;
        RECT 9.400001 15.100000 9.800000 15.200000 ;
        RECT 8.600000 14.800000 9.800000 15.100000 ;
        RECT 13.400001 14.800000 13.800000 15.200000 ;
        RECT 14.200000 14.800000 14.600000 15.200000 ;
        RECT 18.200001 15.100000 18.600000 15.200000 ;
        RECT 19.000000 15.100000 19.400000 15.200000 ;
        RECT 18.200001 14.800000 19.400000 15.100000 ;
        RECT 20.600000 14.200000 20.900000 21.800001 ;
        RECT 1.400000 13.100000 1.800000 13.500000 ;
        RECT 2.100000 13.200000 4.900000 13.500000 ;
        RECT 4.500000 13.100000 4.900000 13.200000 ;
        RECT 9.400001 13.800000 9.800000 14.200000 ;
        RECT 15.800000 14.100000 16.200001 14.200000 ;
        RECT 16.600000 14.100000 17.000000 14.200000 ;
        RECT 15.800000 13.800000 17.000000 14.100000 ;
        RECT 20.600000 13.800000 21.000000 14.200000 ;
        RECT 9.400001 13.200000 9.700000 13.800000 ;
        RECT 20.600000 13.200000 20.900000 13.800000 ;
        RECT 9.400001 12.800000 9.800000 13.200000 ;
        RECT 10.200000 13.100000 10.600000 13.200000 ;
        RECT 11.000000 13.100000 11.400001 13.200000 ;
        RECT 10.200000 12.800000 11.400001 13.100000 ;
        RECT 13.400001 12.800000 13.800000 13.200000 ;
        RECT 20.600000 12.800000 21.000000 13.200000 ;
        RECT 13.400001 12.200000 13.700000 12.800000 ;
        RECT 3.000000 11.800000 3.400000 12.200000 ;
        RECT 10.200000 12.100000 10.600000 12.200000 ;
        RECT 11.000000 12.100000 11.400001 12.200000 ;
        RECT 10.200000 11.800000 11.400001 12.100000 ;
        RECT 13.400001 11.800000 13.800000 12.200000 ;
        RECT 15.000000 11.800000 15.400001 12.200000 ;
        RECT 19.800001 11.800000 20.200001 12.200000 ;
        RECT 3.000000 7.200000 3.300000 11.800000 ;
        RECT 3.800000 7.500000 4.200000 7.900000 ;
        RECT 6.900000 7.800000 7.300000 7.900000 ;
        RECT 4.500000 7.500000 7.300000 7.800000 ;
        RECT 3.000000 6.800000 3.400000 7.200000 ;
        RECT 3.800000 7.100000 4.100000 7.500000 ;
        RECT 4.500000 7.400000 4.900000 7.500000 ;
        RECT 6.200000 7.400000 6.600000 7.500000 ;
        RECT 3.800000 6.800000 6.600000 7.100000 ;
        RECT 3.800000 5.100000 4.100000 6.800000 ;
        RECT 6.300000 6.100000 6.600000 6.800000 ;
        RECT 6.300000 5.700000 6.700000 6.100000 ;
        RECT 7.000000 5.100000 7.300000 7.500000 ;
        RECT 8.600000 7.800000 9.000000 8.200000 ;
        RECT 8.600000 7.200000 8.900001 7.800000 ;
        RECT 7.800000 6.800000 8.200000 7.200000 ;
        RECT 8.600000 6.800000 9.000000 7.200000 ;
        RECT 10.200000 7.100000 10.600000 7.200000 ;
        RECT 11.000000 7.100000 11.400001 7.200000 ;
        RECT 10.200000 6.800000 11.400001 7.100000 ;
        RECT 13.400001 7.100000 13.700000 11.800000 ;
        RECT 14.200000 8.800000 14.600000 9.200000 ;
        RECT 14.200000 8.200000 14.500000 8.800000 ;
        RECT 14.200000 7.800000 14.600000 8.200000 ;
        RECT 14.200000 7.100000 14.600000 7.200000 ;
        RECT 13.400001 6.800000 14.600000 7.100000 ;
        RECT 7.800000 6.200000 8.100000 6.800000 ;
        RECT 7.800000 5.800000 8.200000 6.200000 ;
        RECT 15.000000 6.100000 15.300000 11.800000 ;
        RECT 19.800001 9.200000 20.100000 11.800000 ;
        RECT 21.400000 9.200000 21.700001 25.800001 ;
        RECT 23.100000 25.100000 23.400000 27.500000 ;
        RECT 23.800001 27.400000 24.200001 27.500000 ;
        RECT 25.500000 27.400000 25.900000 27.500000 ;
        RECT 26.300001 27.100000 26.600000 27.500000 ;
        RECT 39.799999 27.200001 40.100002 27.800001 ;
        RECT 44.600002 27.500000 45.000000 27.900000 ;
        RECT 47.700001 27.800001 48.100002 27.900000 ;
        RECT 45.299999 27.500000 48.100002 27.800001 ;
        RECT 23.800001 26.800001 26.600000 27.100000 ;
        RECT 23.800001 26.100000 24.100000 26.800001 ;
        RECT 23.700001 25.700001 24.100000 26.100000 ;
        RECT 26.300001 25.100000 26.600000 26.800001 ;
        RECT 29.400000 26.800001 29.800001 27.200001 ;
        RECT 34.200001 27.100000 34.600002 27.200001 ;
        RECT 35.000000 27.100000 35.400002 27.200001 ;
        RECT 34.200001 26.800001 35.400002 27.100000 ;
        RECT 39.799999 26.800001 40.200001 27.200001 ;
        RECT 44.600002 27.100000 44.900002 27.500000 ;
        RECT 45.299999 27.400000 45.700001 27.500000 ;
        RECT 47.000000 27.400000 47.400002 27.500000 ;
        RECT 44.600002 26.800001 47.400002 27.100000 ;
        RECT 29.400000 26.200001 29.700001 26.800001 ;
        RECT 29.400000 25.800001 29.800001 26.200001 ;
        RECT 33.400002 25.800001 33.799999 26.200001 ;
        RECT 35.799999 25.800001 36.200001 26.200001 ;
        RECT 41.400002 25.800001 41.799999 26.200001 ;
        RECT 23.100000 24.700001 23.500000 25.100000 ;
        RECT 26.200001 24.700001 26.600000 25.100000 ;
        RECT 24.600000 22.100000 25.000000 22.200001 ;
        RECT 25.400000 22.100000 25.800001 22.200001 ;
        RECT 24.600000 21.800001 25.800001 22.100000 ;
        RECT 27.800001 21.800001 28.200001 22.200001 ;
        RECT 30.200001 21.800001 30.600000 22.200001 ;
        RECT 22.200001 16.800001 22.600000 17.200001 ;
        RECT 22.200001 16.200001 22.500000 16.800001 ;
        RECT 22.200001 15.800000 22.600000 16.200001 ;
        RECT 23.000000 15.800000 23.400000 16.200001 ;
        RECT 26.200001 16.100000 26.600000 16.200001 ;
        RECT 27.000000 16.100000 27.400000 16.200001 ;
        RECT 26.200001 15.800000 27.400000 16.100000 ;
        RECT 23.000000 13.200000 23.300001 15.800000 ;
        RECT 27.800001 14.200000 28.100000 21.800001 ;
        RECT 28.600000 15.900001 29.000000 16.300001 ;
        RECT 28.600000 14.200000 28.900000 15.900001 ;
        RECT 30.200001 15.200000 30.500000 21.800001 ;
        RECT 31.700001 15.900001 32.100002 16.300001 ;
        RECT 30.200001 14.800000 30.600000 15.200000 ;
        RECT 31.100000 14.900001 31.500000 15.300000 ;
        RECT 31.100000 14.200000 31.400000 14.900001 ;
        RECT 27.800001 13.800000 28.200001 14.200000 ;
        RECT 28.600000 13.900001 31.400000 14.200000 ;
        RECT 28.600000 13.500000 28.900000 13.900001 ;
        RECT 29.300001 13.500000 29.700001 13.600000 ;
        RECT 31.000000 13.500000 31.400000 13.600000 ;
        RECT 31.800001 13.500000 32.100002 15.900001 ;
        RECT 33.400002 16.200001 33.700001 25.800001 ;
        RECT 35.799999 25.200001 36.100002 25.800001 ;
        RECT 41.400002 25.200001 41.700001 25.800001 ;
        RECT 35.799999 24.800001 36.200001 25.200001 ;
        RECT 38.200001 25.100000 38.600002 25.200001 ;
        RECT 39.000000 25.100000 39.400002 25.200001 ;
        RECT 38.200001 24.800001 39.400002 25.100000 ;
        RECT 41.400002 24.800001 41.799999 25.200001 ;
        RECT 44.600002 25.100000 44.900002 26.800001 ;
        RECT 45.400002 26.100000 45.799999 26.200001 ;
        RECT 46.200001 26.100000 46.600002 26.200001 ;
        RECT 45.400002 25.800001 46.600002 26.100000 ;
        RECT 47.100002 26.100000 47.400002 26.800001 ;
        RECT 47.100002 25.700001 47.500000 26.100000 ;
        RECT 47.799999 25.100000 48.100002 27.500000 ;
        RECT 52.600002 27.500000 53.000000 27.900000 ;
        RECT 55.700001 27.800001 56.100002 27.900000 ;
        RECT 53.299999 27.500000 56.100002 27.800001 ;
        RECT 51.799999 26.800001 52.200001 27.200001 ;
        RECT 52.600002 27.100000 52.900002 27.500000 ;
        RECT 53.299999 27.400000 53.700001 27.500000 ;
        RECT 55.000000 27.400000 55.400002 27.500000 ;
        RECT 52.600002 26.800001 55.400002 27.100000 ;
        RECT 51.799999 26.200001 52.100002 26.800001 ;
        RECT 51.799999 25.800001 52.200001 26.200001 ;
        RECT 44.600002 24.700001 45.000000 25.100000 ;
        RECT 47.700001 24.700001 48.100002 25.100000 ;
        RECT 52.600002 25.100000 52.900002 26.800001 ;
        RECT 53.400002 26.100000 53.799999 26.200001 ;
        RECT 54.200001 26.100000 54.600002 26.200001 ;
        RECT 53.400002 25.800001 54.600002 26.100000 ;
        RECT 55.100002 26.100000 55.400002 26.800001 ;
        RECT 55.100002 25.700001 55.500000 26.100000 ;
        RECT 55.799999 25.100000 56.100002 27.500000 ;
        RECT 52.600002 24.700001 53.000000 25.100000 ;
        RECT 55.700001 24.700001 56.100002 25.100000 ;
        RECT 56.600002 26.800001 57.000000 27.200001 ;
        RECT 39.799999 23.800001 40.200001 24.200001 ;
        RECT 35.799999 21.800001 36.200001 22.200001 ;
        RECT 33.400002 15.800000 33.799999 16.200001 ;
        RECT 33.400002 14.200000 33.700001 15.800000 ;
        RECT 35.799999 14.200000 36.100002 21.800001 ;
        RECT 39.000000 15.800000 39.400002 16.200001 ;
        RECT 39.799999 16.100000 40.100002 23.800001 ;
        RECT 56.600002 19.200001 56.900002 26.800001 ;
        RECT 58.200001 25.800001 58.600002 26.200001 ;
        RECT 61.400002 25.800001 61.799999 26.200001 ;
        RECT 58.200001 25.200001 58.500000 25.800001 ;
        RECT 58.200001 24.800001 58.600002 25.200001 ;
        RECT 57.400002 21.800001 57.799999 22.200001 ;
        RECT 53.400002 18.800001 53.799999 19.200001 ;
        RECT 56.600002 18.800001 57.000000 19.200001 ;
        RECT 42.200001 17.100000 42.600002 17.200001 ;
        RECT 43.000000 17.100000 43.400002 17.200001 ;
        RECT 42.200001 16.800001 43.400002 17.100000 ;
        RECT 45.400002 16.800001 45.799999 17.200001 ;
        RECT 45.400002 16.200001 45.700001 16.800001 ;
        RECT 40.600002 16.100000 41.000000 16.200001 ;
        RECT 39.799999 15.800000 41.000000 16.100000 ;
        RECT 42.200001 16.100000 42.600002 16.200001 ;
        RECT 43.000000 16.100000 43.400002 16.200001 ;
        RECT 42.200001 15.800000 43.400002 16.100000 ;
        RECT 45.400002 15.800000 45.799999 16.200001 ;
        RECT 39.000000 15.200000 39.299999 15.800000 ;
        RECT 40.600002 15.200000 40.900002 15.800000 ;
        RECT 39.000000 14.800000 39.400002 15.200000 ;
        RECT 40.600002 14.800000 41.000000 15.200000 ;
        RECT 43.000000 14.800000 43.400002 15.200000 ;
        RECT 43.000000 14.200000 43.299999 14.800000 ;
        RECT 53.400002 14.200000 53.700001 18.800001 ;
        RECT 57.400002 17.200001 57.700001 21.800001 ;
        RECT 57.400002 16.800001 57.799999 17.200001 ;
        RECT 54.200001 15.800000 54.600002 16.200001 ;
        RECT 57.400002 15.900001 57.799999 16.300001 ;
        RECT 59.000000 16.100000 59.400002 16.200001 ;
        RECT 59.799999 16.100000 60.200001 16.200001 ;
        RECT 23.000000 12.800000 23.400000 13.200000 ;
        RECT 23.800001 12.800000 24.200001 13.200000 ;
        RECT 28.600000 13.100000 29.000000 13.500000 ;
        RECT 29.300001 13.200000 32.100002 13.500000 ;
        RECT 31.700001 13.100000 32.100002 13.200000 ;
        RECT 32.600002 13.800000 33.000000 14.200000 ;
        RECT 33.400002 13.800000 33.799999 14.200000 ;
        RECT 35.799999 13.800000 36.200001 14.200000 ;
        RECT 39.000000 14.100000 39.400002 14.200000 ;
        RECT 39.799999 14.100000 40.200001 14.200000 ;
        RECT 39.000000 13.800000 40.200001 14.100000 ;
        RECT 43.000000 13.800000 43.400002 14.200000 ;
        RECT 44.600002 14.100000 45.000000 14.200000 ;
        RECT 45.400002 14.100000 45.799999 14.200000 ;
        RECT 44.600002 13.800000 45.799999 14.100000 ;
        RECT 47.000000 14.100000 47.400002 14.200000 ;
        RECT 47.799999 14.100000 48.200001 14.200000 ;
        RECT 47.000000 13.800000 48.200001 14.100000 ;
        RECT 52.600002 14.100000 53.000000 14.200000 ;
        RECT 53.400002 14.100000 53.799999 14.200000 ;
        RECT 52.600002 13.800000 53.799999 14.100000 ;
        RECT 32.600002 13.200000 32.900002 13.800000 ;
        RECT 35.799999 13.200000 36.100002 13.800000 ;
        RECT 54.200001 13.200000 54.500000 15.800000 ;
        RECT 57.400002 14.200000 57.700001 15.900001 ;
        RECT 59.000000 15.800000 60.200001 16.100000 ;
        RECT 60.500000 15.900001 60.900002 16.300001 ;
        RECT 59.900002 14.900001 60.299999 15.300000 ;
        RECT 59.900002 14.200000 60.200001 14.900001 ;
        RECT 55.799999 13.800000 56.200001 14.200000 ;
        RECT 56.600002 13.800000 57.000000 14.200000 ;
        RECT 57.400002 13.900001 60.200001 14.200000 ;
        RECT 32.600002 12.800000 33.000000 13.200000 ;
        RECT 35.799999 12.800000 36.200001 13.200000 ;
        RECT 38.200001 13.100000 38.600002 13.200000 ;
        RECT 39.000000 13.100000 39.400002 13.200000 ;
        RECT 38.200001 12.800000 39.400002 13.100000 ;
        RECT 43.000000 12.800000 43.400002 13.200000 ;
        RECT 50.200001 12.800000 50.600002 13.200000 ;
        RECT 54.200001 12.800000 54.600002 13.200000 ;
        RECT 23.800001 12.200000 24.100000 12.800000 ;
        RECT 23.800001 11.800000 24.200001 12.200000 ;
        RECT 26.200001 11.800000 26.600000 12.200000 ;
        RECT 30.200001 11.800000 30.600000 12.200000 ;
        RECT 33.400002 11.800000 33.799999 12.200000 ;
        RECT 36.600002 11.800000 37.000000 12.200000 ;
        RECT 19.800001 8.800000 20.200001 9.200000 ;
        RECT 21.400000 8.800000 21.800001 9.200000 ;
        RECT 22.200001 9.100000 22.600000 9.200000 ;
        RECT 23.000000 9.100000 23.400000 9.200000 ;
        RECT 22.200001 8.800000 23.400000 9.100000 ;
        RECT 26.200001 8.200000 26.500000 11.800000 ;
        RECT 29.400000 8.800000 29.800001 9.200000 ;
        RECT 29.400000 8.200000 29.700001 8.800000 ;
        RECT 22.200001 7.800000 22.600000 8.200000 ;
        RECT 26.200001 7.800000 26.600000 8.200000 ;
        RECT 29.400000 7.800000 29.800001 8.200000 ;
        RECT 22.200001 7.200000 22.500000 7.800000 ;
        RECT 22.200001 7.100000 22.600000 7.200000 ;
        RECT 23.000000 7.100000 23.400000 7.200000 ;
        RECT 30.200001 7.100000 30.500000 11.800000 ;
        RECT 22.200001 6.800000 23.400000 7.100000 ;
        RECT 29.400000 6.800000 30.500000 7.100000 ;
        RECT 29.400000 6.200000 29.700001 6.800000 ;
        RECT 15.800000 6.100000 16.200001 6.200000 ;
        RECT 15.000000 5.800000 16.200001 6.100000 ;
        RECT 29.400000 5.800000 29.800001 6.200000 ;
        RECT 15.000000 5.200000 15.300000 5.800000 ;
        RECT 33.400002 5.200000 33.700001 11.800000 ;
        RECT 35.799999 7.800000 36.200001 8.200000 ;
        RECT 35.799999 7.200000 36.100002 7.800000 ;
        RECT 35.799999 6.800000 36.200001 7.200000 ;
        RECT 36.600002 5.200000 36.900002 11.800000 ;
        RECT 43.000000 9.200000 43.299999 12.800000 ;
        RECT 45.400002 12.100000 45.799999 12.200000 ;
        RECT 46.200001 12.100000 46.600002 12.200000 ;
        RECT 45.400002 11.800000 46.600002 12.100000 ;
        RECT 50.200001 9.200000 50.500000 12.800000 ;
        RECT 51.000000 11.800000 51.400002 12.200000 ;
        RECT 51.000000 9.200000 51.299999 11.800000 ;
        RECT 55.799999 9.200000 56.100002 13.800000 ;
        RECT 56.600002 12.200000 56.900002 13.800000 ;
        RECT 57.400002 13.500000 57.700001 13.900001 ;
        RECT 58.100002 13.500000 58.500000 13.600000 ;
        RECT 59.799999 13.500000 60.200001 13.600000 ;
        RECT 60.600002 13.500000 60.900002 15.900001 ;
        RECT 61.400002 15.200000 61.700001 25.800001 ;
        RECT 62.200001 15.800000 62.600002 16.200001 ;
        RECT 62.200001 15.200000 62.500000 15.800000 ;
        RECT 61.400002 14.800000 61.799999 15.200000 ;
        RECT 62.200001 14.800000 62.600002 15.200000 ;
        RECT 57.400002 13.100000 57.799999 13.500000 ;
        RECT 58.100002 13.200000 60.900002 13.500000 ;
        RECT 60.500000 13.100000 60.900002 13.200000 ;
        RECT 61.400002 13.800000 61.799999 14.200000 ;
        RECT 61.400002 13.200000 61.700001 13.800000 ;
        RECT 61.400002 12.800000 61.799999 13.200000 ;
        RECT 56.600002 11.800000 57.000000 12.200000 ;
        RECT 39.799999 9.100000 40.200001 9.200000 ;
        RECT 40.600002 9.100000 41.000000 9.200000 ;
        RECT 39.799999 8.800000 41.000000 9.100000 ;
        RECT 43.000000 8.800000 43.400002 9.200000 ;
        RECT 50.200001 8.800000 50.600002 9.200000 ;
        RECT 51.000000 8.800000 51.400002 9.200000 ;
        RECT 55.799999 8.800000 56.200001 9.200000 ;
        RECT 59.799999 9.100000 60.200001 9.200000 ;
        RECT 60.600002 9.100000 61.000000 9.200000 ;
        RECT 59.799999 8.800000 61.000000 9.100000 ;
        RECT 48.600002 7.500000 49.000000 7.900000 ;
        RECT 51.700001 7.800000 52.100002 7.900000 ;
        RECT 49.299999 7.500000 52.100002 7.800000 ;
        RECT 39.000000 6.800000 39.400002 7.200000 ;
        RECT 40.600002 7.100000 41.000000 7.200000 ;
        RECT 41.400002 7.100000 41.799999 7.200000 ;
        RECT 40.600002 6.800000 41.799999 7.100000 ;
        RECT 43.000000 6.800000 43.400002 7.200000 ;
        RECT 48.600002 7.100000 48.900002 7.500000 ;
        RECT 49.299999 7.400000 49.700001 7.500000 ;
        RECT 51.000000 7.400000 51.400002 7.500000 ;
        RECT 48.600002 6.800000 51.400002 7.100000 ;
        RECT 39.000000 6.200000 39.299999 6.800000 ;
        RECT 43.000000 6.200000 43.299999 6.800000 ;
        RECT 39.000000 5.800000 39.400002 6.200000 ;
        RECT 40.600002 6.100000 41.000000 6.200000 ;
        RECT 41.400002 6.100000 41.799999 6.200000 ;
        RECT 40.600002 5.800000 41.799999 6.100000 ;
        RECT 43.000000 5.800000 43.400002 6.200000 ;
        RECT 3.800000 4.700000 4.200000 5.100000 ;
        RECT 6.900000 4.700000 7.300000 5.100000 ;
        RECT 10.200000 5.100000 10.600000 5.200000 ;
        RECT 11.000000 5.100000 11.400001 5.200000 ;
        RECT 10.200000 4.800000 11.400001 5.100000 ;
        RECT 15.000000 4.800000 15.400001 5.200000 ;
        RECT 33.400002 4.800000 33.799999 5.200000 ;
        RECT 36.600002 4.800000 37.000000 5.200000 ;
        RECT 48.600002 5.100000 48.900002 6.800000 ;
        RECT 51.100002 6.100000 51.400002 6.800000 ;
        RECT 51.100002 5.700000 51.500000 6.100000 ;
        RECT 51.799999 5.100000 52.100002 7.500000 ;
        RECT 58.299999 7.800000 58.700001 7.900000 ;
        RECT 58.299999 7.500000 61.100002 7.800000 ;
        RECT 61.400002 7.500000 61.799999 7.900000 ;
        RECT 55.799999 6.100000 56.200001 6.200000 ;
        RECT 56.600002 6.100000 57.000000 6.200000 ;
        RECT 55.799999 5.800000 57.000000 6.100000 ;
        RECT 48.600002 4.700000 49.000000 5.100000 ;
        RECT 51.700001 4.700000 52.100002 5.100000 ;
        RECT 58.299999 5.100000 58.600002 7.500000 ;
        RECT 59.000000 7.400000 59.400002 7.500000 ;
        RECT 60.700001 7.400000 61.100002 7.500000 ;
        RECT 61.500000 7.100000 61.799999 7.500000 ;
        RECT 59.000000 6.800000 61.799999 7.100000 ;
        RECT 59.000000 6.100000 59.299999 6.800000 ;
        RECT 58.900002 5.700000 59.299999 6.100000 ;
        RECT 61.500000 5.100000 61.799999 6.800000 ;
        RECT 58.299999 4.700000 58.700001 5.100000 ;
        RECT 61.400002 4.700000 61.799999 5.100000 ;
      LAYER via2 ;
        RECT 11.000000 28.800001 11.400001 29.200001 ;
        RECT 38.200001 27.800001 38.600002 28.200001 ;
        RECT 19.000000 21.800001 19.400000 22.200001 ;
        RECT 16.600000 13.800000 17.000000 14.200000 ;
        RECT 11.000000 11.800000 11.400001 12.200000 ;
        RECT 39.000000 24.800001 39.400002 25.200001 ;
        RECT 46.200001 25.800001 46.600002 26.200001 ;
        RECT 43.000000 16.800001 43.400002 17.200001 ;
        RECT 40.600002 15.800000 41.000000 16.200001 ;
        RECT 45.400002 13.800000 45.799999 14.200000 ;
        RECT 47.799999 13.800000 48.200001 14.200000 ;
        RECT 59.799999 15.800000 60.200001 16.200001 ;
        RECT 39.000000 12.800000 39.400002 13.200000 ;
        RECT 23.000000 6.800000 23.400000 7.200000 ;
        RECT 46.200001 11.800000 46.600002 12.200000 ;
        RECT 40.600002 8.800000 41.000000 9.200000 ;
        RECT 60.600002 8.800000 61.000000 9.200000 ;
        RECT 41.400002 5.800000 41.799999 6.200000 ;
        RECT 11.000000 4.800000 11.400001 5.200000 ;
      LAYER metal3 ;
        RECT 7.800000 29.100000 8.200000 29.200001 ;
        RECT 11.000000 29.100000 11.400001 29.200001 ;
        RECT 7.800000 28.800001 11.400001 29.100000 ;
        RECT 38.200001 28.100000 38.600002 28.200001 ;
        RECT 39.799999 28.100000 40.200001 28.200001 ;
        RECT 38.200001 27.800001 40.200001 28.100000 ;
        RECT 29.400000 27.100000 29.800001 27.200001 ;
        RECT 34.200001 27.100000 34.600002 27.200001 ;
        RECT 29.400000 26.800001 34.600002 27.100000 ;
        RECT 1.400000 26.100000 1.800000 26.200001 ;
        RECT 46.200001 26.100000 46.600002 26.200001 ;
        RECT 51.799999 26.100000 52.200001 26.200001 ;
        RECT 1.400000 25.800001 5.700000 26.100000 ;
        RECT 46.200001 25.800001 52.200001 26.100000 ;
        RECT 53.400002 26.100000 53.799999 26.200001 ;
        RECT 58.200001 26.100000 58.600002 26.200001 ;
        RECT 53.400002 25.800001 58.600002 26.100000 ;
        RECT 5.400000 25.200001 5.700000 25.800001 ;
        RECT 3.000000 25.100000 3.400000 25.200001 ;
        RECT 3.800000 25.100000 4.200000 25.200001 ;
        RECT 3.000000 24.800001 4.200000 25.100000 ;
        RECT 5.400000 24.800001 5.800000 25.200001 ;
        RECT 35.799999 25.100000 36.200001 25.200001 ;
        RECT 39.000000 25.100000 39.400002 25.200001 ;
        RECT 41.400002 25.100000 41.799999 25.200001 ;
        RECT 35.799999 24.800001 41.799999 25.100000 ;
        RECT 19.000000 22.100000 19.400000 22.200001 ;
        RECT 20.600000 22.100000 21.000000 22.200001 ;
        RECT 19.000000 21.800001 21.000000 22.100000 ;
        RECT 24.600000 22.100000 25.000000 22.200001 ;
        RECT 27.800001 22.100000 28.200001 22.200001 ;
        RECT 24.600000 21.800001 28.200001 22.100000 ;
        RECT 53.400002 19.100000 53.799999 19.200001 ;
        RECT 56.600002 19.100000 57.000000 19.200001 ;
        RECT 53.400002 18.800001 57.000000 19.100000 ;
        RECT 22.200001 16.800001 22.600000 17.200001 ;
        RECT 43.000000 17.100000 43.400002 17.200001 ;
        RECT 45.400002 17.100000 45.799999 17.200001 ;
        RECT 42.200001 16.800001 45.799999 17.100000 ;
        RECT 56.600002 17.100000 57.000000 17.200001 ;
        RECT 57.400002 17.100000 57.799999 17.200001 ;
        RECT 56.600002 16.800001 57.799999 17.100000 ;
        RECT 22.200001 16.100000 22.500000 16.800001 ;
        RECT 26.200001 16.100000 26.600000 16.200001 ;
        RECT 22.200001 15.800000 26.600000 16.100000 ;
        RECT 40.600002 16.100000 41.000000 16.200001 ;
        RECT 42.200001 16.100000 42.600002 16.200001 ;
        RECT 40.600002 15.800000 42.600002 16.100000 ;
        RECT 59.799999 16.100000 60.200001 16.200001 ;
        RECT 62.200001 16.100000 62.600002 16.200001 ;
        RECT 59.799999 15.800000 62.600002 16.100000 ;
        RECT 7.800000 15.100000 8.200000 15.200000 ;
        RECT 8.600000 15.100000 9.000000 15.200000 ;
        RECT 13.400001 15.100000 13.800000 15.200000 ;
        RECT 7.800000 14.800000 13.800000 15.100000 ;
        RECT 14.200000 15.100000 14.600000 15.200000 ;
        RECT 18.200001 15.100000 18.600000 15.200000 ;
        RECT 14.200000 14.800000 18.600000 15.100000 ;
        RECT 29.400000 15.100000 29.800001 15.200000 ;
        RECT 30.200001 15.100000 30.600000 15.200000 ;
        RECT 29.400000 14.800000 30.600000 15.100000 ;
        RECT 39.000000 15.100000 39.400002 15.200000 ;
        RECT 43.000000 15.100000 43.400002 15.200000 ;
        RECT 39.000000 14.800000 43.400002 15.100000 ;
        RECT 59.799999 15.100000 60.200001 15.200000 ;
        RECT 61.400002 15.100000 61.799999 15.200000 ;
        RECT 59.799999 14.800000 61.799999 15.100000 ;
        RECT 16.600000 14.100000 17.000000 14.200000 ;
        RECT 20.600000 14.100000 21.000000 14.200000 ;
        RECT 16.600000 13.800000 21.000000 14.100000 ;
        RECT 33.400002 14.100000 33.799999 14.200000 ;
        RECT 39.000000 14.100000 39.400002 14.200000 ;
        RECT 33.400002 13.800000 39.400002 14.100000 ;
        RECT 45.400002 14.100000 45.799999 14.200000 ;
        RECT 47.799999 14.100000 48.200001 14.200000 ;
        RECT 52.600002 14.100000 53.000000 14.200000 ;
        RECT 45.400002 13.800000 53.000000 14.100000 ;
        RECT 55.799999 14.100000 56.200001 14.200000 ;
        RECT 55.799999 13.800000 61.700001 14.100000 ;
        RECT 61.400002 13.200000 61.700001 13.800000 ;
        RECT 9.400001 13.100000 9.800000 13.200000 ;
        RECT 10.200000 13.100000 10.600000 13.200000 ;
        RECT 9.400001 12.800000 10.600000 13.100000 ;
        RECT 13.400001 13.100000 13.800000 13.200000 ;
        RECT 23.000000 13.100000 23.400000 13.200000 ;
        RECT 13.400001 12.800000 23.400000 13.100000 ;
        RECT 32.600002 13.100000 33.000000 13.200000 ;
        RECT 39.000000 13.100000 39.400002 13.200000 ;
        RECT 32.600002 12.800000 39.400002 13.100000 ;
        RECT 43.000000 13.100000 43.400002 13.200000 ;
        RECT 54.200001 13.100000 54.600002 13.200000 ;
        RECT 43.000000 12.800000 54.600002 13.100000 ;
        RECT 61.400002 12.800000 61.799999 13.200000 ;
        RECT 11.000000 12.100000 11.400001 12.200000 ;
        RECT 23.800001 12.100000 24.200001 12.200000 ;
        RECT 10.200000 11.800000 24.200001 12.100000 ;
        RECT 36.600002 12.100000 37.000000 12.200000 ;
        RECT 46.200001 12.100000 46.600002 12.200000 ;
        RECT 36.600002 11.800000 46.600002 12.100000 ;
        RECT 51.000000 12.100000 51.400002 12.200000 ;
        RECT 56.600002 12.100000 57.000000 12.200000 ;
        RECT 51.000000 11.800000 57.000000 12.100000 ;
        RECT 14.200000 9.100000 14.600000 9.200000 ;
        RECT 19.800001 9.100000 20.200001 9.200000 ;
        RECT 14.200000 8.800000 20.200001 9.100000 ;
        RECT 21.400000 9.100000 21.800001 9.200000 ;
        RECT 22.200001 9.100000 22.600000 9.200000 ;
        RECT 21.400000 8.800000 22.600000 9.100000 ;
        RECT 29.400000 8.800000 29.800001 9.200000 ;
        RECT 40.600002 9.100000 41.000000 9.200000 ;
        RECT 50.200001 9.100000 50.600002 9.200000 ;
        RECT 39.799999 8.800000 50.600002 9.100000 ;
        RECT 59.799999 9.100000 60.200001 9.200000 ;
        RECT 60.600002 9.100000 61.000000 9.200000 ;
        RECT 59.799999 8.800000 61.000000 9.100000 ;
        RECT 29.400000 8.200000 29.700001 8.800000 ;
        RECT 3.000000 8.100000 3.400000 8.200000 ;
        RECT 8.600000 8.100000 9.000000 8.200000 ;
        RECT 22.200001 8.100000 22.600000 8.200000 ;
        RECT 3.000000 7.800000 22.600000 8.100000 ;
        RECT 29.400000 7.800000 29.800001 8.200000 ;
        RECT 35.799999 7.800000 36.200001 8.200000 ;
        RECT 10.200000 7.100000 10.600000 7.200000 ;
        RECT 7.800000 6.800000 10.600000 7.100000 ;
        RECT 23.000000 7.100000 23.400000 7.200000 ;
        RECT 35.799999 7.100000 36.100002 7.800000 ;
        RECT 23.000000 6.800000 36.100002 7.100000 ;
        RECT 39.000000 7.100000 39.400002 7.200000 ;
        RECT 40.600002 7.100000 41.000000 7.200000 ;
        RECT 39.000000 6.800000 41.000000 7.100000 ;
        RECT 7.800000 6.200000 8.100000 6.800000 ;
        RECT 7.800000 5.800000 8.200000 6.200000 ;
        RECT 41.400002 6.100000 41.799999 6.200000 ;
        RECT 43.000000 6.100000 43.400002 6.200000 ;
        RECT 41.400002 5.800000 43.400002 6.100000 ;
        RECT 55.799999 6.100000 56.200001 6.200000 ;
        RECT 56.600002 6.100000 57.000000 6.200000 ;
        RECT 55.799999 5.800000 57.000000 6.100000 ;
        RECT 11.000000 5.100000 11.400001 5.200000 ;
        RECT 15.000000 5.100000 15.400001 5.200000 ;
        RECT 11.000000 4.800000 15.400001 5.100000 ;
      LAYER via3 ;
        RECT 3.800000 24.800001 4.200000 25.200001 ;
        RECT 56.600002 5.800000 57.000000 6.200000 ;
      LAYER metal4 ;
        RECT 3.800000 25.100000 4.200000 25.200001 ;
        RECT 3.000000 24.800001 4.200000 25.100000 ;
        RECT 3.000000 8.200000 3.300000 24.800001 ;
        RECT 56.600002 16.800001 57.000000 17.200001 ;
        RECT 29.400000 14.800000 29.800001 15.200000 ;
        RECT 29.400000 8.200000 29.700001 14.800000 ;
        RECT 3.000000 7.800000 3.400000 8.200000 ;
        RECT 29.400000 7.800000 29.800001 8.200000 ;
        RECT 56.600002 6.200000 56.900002 16.800001 ;
        RECT 59.799999 14.800000 60.200001 15.200000 ;
        RECT 59.799999 9.200000 60.100002 14.800000 ;
        RECT 59.799999 8.800000 60.200001 9.200000 ;
        RECT 56.600002 5.800000 57.000000 6.200000 ;
  END
END adder
