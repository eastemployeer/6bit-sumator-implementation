magic
tech scmos
magscale 1 2
timestamp 1591288394
<< metal1 >>
rect 314 214 326 216
rect 299 206 301 214
rect 309 206 311 214
rect 319 206 321 214
rect 329 206 331 214
rect 339 206 341 214
rect 314 204 326 206
rect 125 157 204 163
rect 292 137 371 143
rect 461 137 476 143
rect 93 117 115 123
rect 132 117 227 123
rect 285 117 300 123
rect 420 117 435 123
rect 138 14 150 16
rect 123 6 125 14
rect 133 6 135 14
rect 143 6 145 14
rect 153 6 155 14
rect 163 6 165 14
rect 138 4 150 6
<< m2contact >>
rect 291 206 299 214
rect 301 206 309 214
rect 311 206 319 214
rect 321 206 329 214
rect 331 206 339 214
rect 341 206 349 214
rect 12 156 20 164
rect 204 156 212 164
rect 252 156 260 164
rect 268 156 276 164
rect 60 136 68 144
rect 284 136 292 144
rect 476 136 484 144
rect 44 116 52 124
rect 124 116 132 124
rect 236 116 244 124
rect 300 116 308 124
rect 380 116 388 124
rect 412 116 420 124
rect 115 6 123 14
rect 125 6 133 14
rect 135 6 143 14
rect 145 6 153 14
rect 155 6 163 14
rect 165 6 173 14
<< metal2 >>
rect 253 184 259 263
rect 314 214 326 216
rect 299 206 301 214
rect 309 206 311 214
rect 319 206 321 214
rect 329 206 331 214
rect 339 206 341 214
rect 314 204 326 206
rect 253 164 259 176
rect 285 144 291 176
rect 301 124 307 156
rect 381 124 387 156
rect 477 124 483 136
rect 138 14 150 16
rect 123 6 125 14
rect 133 6 135 14
rect 143 6 145 14
rect 153 6 155 14
rect 163 6 165 14
rect 138 4 150 6
<< m3contact >>
rect 291 206 299 214
rect 301 206 309 214
rect 311 206 319 214
rect 321 206 329 214
rect 331 206 339 214
rect 341 206 349 214
rect 252 176 260 184
rect 284 176 292 184
rect 12 156 20 164
rect 204 156 212 164
rect 268 156 276 164
rect 300 156 308 164
rect 380 156 388 164
rect 60 136 68 144
rect 44 116 52 124
rect 124 116 132 124
rect 236 116 244 124
rect 412 116 420 124
rect 476 116 484 124
rect 115 6 123 14
rect 125 6 133 14
rect 135 6 143 14
rect 145 6 153 14
rect 155 6 163 14
rect 165 6 173 14
<< metal3 >>
rect 290 214 350 216
rect 290 206 291 214
rect 300 206 301 214
rect 339 206 340 214
rect 349 206 350 214
rect 290 204 350 206
rect 260 177 284 183
rect -35 157 12 163
rect 212 157 268 163
rect 308 157 380 163
rect 388 157 515 163
rect -35 137 60 143
rect -35 117 -29 137
rect 52 117 124 123
rect 244 117 412 123
rect 484 117 515 123
rect 114 14 174 16
rect 114 6 115 14
rect 124 6 125 14
rect 163 6 164 14
rect 173 6 174 14
rect 114 4 174 6
<< m4contact >>
rect 292 206 299 214
rect 299 206 300 214
rect 304 206 309 214
rect 309 206 311 214
rect 311 206 312 214
rect 316 206 319 214
rect 319 206 321 214
rect 321 206 324 214
rect 328 206 329 214
rect 329 206 331 214
rect 331 206 336 214
rect 340 206 341 214
rect 341 206 348 214
rect 116 6 123 14
rect 123 6 124 14
rect 128 6 133 14
rect 133 6 135 14
rect 135 6 136 14
rect 140 6 143 14
rect 143 6 145 14
rect 145 6 148 14
rect 152 6 153 14
rect 153 6 155 14
rect 155 6 160 14
rect 164 6 165 14
rect 165 6 172 14
<< metal4 >>
rect 112 14 176 216
rect 112 6 116 14
rect 124 6 128 14
rect 136 6 140 14
rect 148 6 152 14
rect 160 6 164 14
rect 172 6 176 14
rect 112 -10 176 6
rect 288 214 352 216
rect 288 206 292 214
rect 300 206 304 214
rect 312 206 316 214
rect 324 206 328 214
rect 336 206 340 214
rect 348 206 352 214
rect 288 -10 352 206
use BUFX2  _9_
timestamp 1591288394
transform -1 0 56 0 -1 210
box -4 -6 52 206
use BUFX2  _10_
timestamp 1591288394
transform -1 0 104 0 -1 210
box -4 -6 52 206
use INVX1  _6_
timestamp 1591288394
transform -1 0 136 0 -1 210
box -4 -6 36 206
use FILL  SFILL1360x100
timestamp 1591288394
transform -1 0 152 0 -1 210
box -4 -6 20 206
use FILL  SFILL1520x100
timestamp 1591288394
transform -1 0 168 0 -1 210
box -4 -6 20 206
use NOR2X1  _7_
timestamp 1591288394
transform 1 0 200 0 -1 210
box -4 -6 52 206
use FILL  SFILL1680x100
timestamp 1591288394
transform -1 0 184 0 -1 210
box -4 -6 20 206
use FILL  SFILL1840x100
timestamp 1591288394
transform -1 0 200 0 -1 210
box -4 -6 20 206
use NOR2X1  _5_
timestamp 1591288394
transform 1 0 248 0 -1 210
box -4 -6 52 206
use FILL  SFILL2960x100
timestamp 1591288394
transform -1 0 312 0 -1 210
box -4 -6 20 206
use AND2X2  _4_
timestamp 1591288394
transform 1 0 360 0 -1 210
box -4 -6 68 206
use FILL  SFILL3120x100
timestamp 1591288394
transform -1 0 328 0 -1 210
box -4 -6 20 206
use FILL  SFILL3280x100
timestamp 1591288394
transform -1 0 344 0 -1 210
box -4 -6 20 206
use FILL  SFILL3440x100
timestamp 1591288394
transform -1 0 360 0 -1 210
box -4 -6 20 206
use BUFX2  _8_
timestamp 1591288394
transform 1 0 424 0 -1 210
box -4 -6 52 206
<< labels >>
flabel metal4 s 112 -10 176 0 7 FreeSans 24 270 0 0 vdd
port 0 nsew default bidirectional
flabel metal4 s 288 -10 352 0 7 FreeSans 24 270 0 0 gnd
port 1 nsew default bidirectional
flabel metal3 s 509 117 515 123 3 FreeSans 24 0 0 0 g
port 2 nsew default bidirectional
flabel metal3 s -35 157 -29 163 7 FreeSans 24 0 0 0 h
port 3 nsew default bidirectional
flabel metal3 s -35 117 -29 123 7 FreeSans 24 0 0 0 p
port 4 nsew default bidirectional
flabel metal3 s 509 157 515 163 3 FreeSans 24 0 0 0 x
port 5 nsew default bidirectional
flabel metal2 s 253 257 259 263 3 FreeSans 24 90 0 0 y
port 6 nsew default bidirectional
<< end >>
