magic
tech scmos
timestamp 1592523827
<< metal1 >>
rect 469 307 475 308
rect 464 303 465 307
rect 469 303 470 307
rect 474 303 475 307
rect 479 303 480 307
rect 469 302 475 303
rect 106 288 108 292
rect 286 278 297 281
rect 142 271 145 278
rect 134 268 145 271
rect 286 268 297 271
rect 430 271 433 281
rect 402 268 409 271
rect 430 268 438 271
rect 294 262 297 268
rect 310 258 329 261
rect 338 258 345 261
rect 458 258 465 261
rect 582 258 593 261
rect 326 248 337 251
rect 414 251 417 258
rect 582 252 585 258
rect 414 248 425 251
rect 146 238 153 241
rect 390 238 398 241
rect 630 238 646 241
rect 166 218 182 221
rect 250 218 254 222
rect 306 218 307 222
rect 173 207 179 208
rect 168 203 169 207
rect 173 203 174 207
rect 178 203 179 207
rect 183 203 184 207
rect 173 202 179 203
rect 78 151 81 158
rect 70 148 81 151
rect 534 151 537 161
rect 430 148 441 151
rect 534 148 553 151
rect 430 142 433 148
rect 110 138 121 141
rect 198 138 217 141
rect 246 138 257 141
rect 350 138 358 141
rect 366 138 377 141
rect 510 138 521 141
rect 526 138 534 141
rect 638 138 646 141
rect 94 131 97 138
rect 86 128 97 131
rect 110 132 113 138
rect 149 118 150 122
rect 266 118 267 122
rect 469 107 475 108
rect 464 103 465 107
rect 469 103 470 107
rect 474 103 475 107
rect 479 103 480 107
rect 469 102 475 103
rect 508 88 510 92
rect 322 78 337 81
rect 114 68 121 71
rect 126 68 137 71
rect 146 68 153 71
rect 246 68 257 71
rect 302 68 313 71
rect 342 68 353 71
rect 390 71 393 81
rect 446 78 473 81
rect 374 68 393 71
rect 470 71 473 78
rect 470 68 481 71
rect 550 71 553 81
rect 534 68 553 71
rect 622 68 630 71
rect 390 62 393 68
rect 22 58 57 61
rect 94 58 113 61
rect 286 58 294 61
rect 430 61 433 68
rect 478 61 481 68
rect 430 58 441 61
rect 478 58 494 61
rect 110 48 113 58
rect 174 48 209 51
rect 214 48 233 51
rect 326 48 334 51
rect 430 48 441 51
rect 173 7 179 8
rect 168 3 169 7
rect 173 3 174 7
rect 178 3 179 7
rect 183 3 184 7
rect 173 2 179 3
<< m2contact >>
rect 460 303 464 307
rect 465 303 469 307
rect 470 303 474 307
rect 475 303 479 307
rect 480 303 484 307
rect 102 288 106 292
rect 198 288 202 292
rect 606 288 610 292
rect 142 278 146 282
rect 158 278 162 282
rect 278 278 282 282
rect 318 278 322 282
rect 374 278 378 282
rect 414 278 418 282
rect 30 268 34 272
rect 78 268 82 272
rect 86 268 90 272
rect 222 268 226 272
rect 270 268 274 272
rect 350 268 354 272
rect 398 268 402 272
rect 582 278 586 282
rect 438 268 442 272
rect 486 268 490 272
rect 518 268 522 272
rect 566 268 570 272
rect 22 258 26 262
rect 54 258 58 262
rect 214 258 218 262
rect 294 258 298 262
rect 334 258 338 262
rect 358 258 362 262
rect 414 258 418 262
rect 454 258 458 262
rect 542 258 546 262
rect 614 258 618 262
rect 382 248 386 252
rect 582 248 586 252
rect 6 238 10 242
rect 142 238 146 242
rect 398 238 402 242
rect 646 238 650 242
rect 182 218 186 222
rect 254 218 258 222
rect 302 218 306 222
rect 358 218 362 222
rect 574 218 578 222
rect 164 203 168 207
rect 169 203 173 207
rect 174 203 178 207
rect 179 203 183 207
rect 184 203 188 207
rect 422 168 426 172
rect 78 158 82 162
rect 134 158 138 162
rect 142 158 146 162
rect 222 158 226 162
rect 230 158 234 162
rect 270 158 274 162
rect 334 158 338 162
rect 390 158 394 162
rect 430 158 434 162
rect 454 158 458 162
rect 94 148 98 152
rect 190 148 194 152
rect 406 148 410 152
rect 542 158 546 162
rect 590 158 594 162
rect 622 148 626 152
rect 6 138 10 142
rect 54 138 58 142
rect 94 138 98 142
rect 158 138 162 142
rect 278 138 282 142
rect 326 138 330 142
rect 358 138 362 142
rect 398 138 402 142
rect 430 138 434 142
rect 446 138 450 142
rect 470 138 474 142
rect 534 138 538 142
rect 558 138 562 142
rect 566 138 570 142
rect 614 138 618 142
rect 646 138 650 142
rect 62 128 66 132
rect 78 128 82 132
rect 110 128 114 132
rect 206 128 210 132
rect 238 128 242 132
rect 358 128 362 132
rect 382 128 386 132
rect 502 128 506 132
rect 30 118 34 122
rect 102 118 106 122
rect 134 118 138 122
rect 150 118 154 122
rect 198 118 202 122
rect 262 118 266 122
rect 302 118 306 122
rect 334 118 338 122
rect 454 118 458 122
rect 460 103 464 107
rect 465 103 469 107
rect 470 103 474 107
rect 475 103 479 107
rect 480 103 484 107
rect 230 88 234 92
rect 398 88 402 92
rect 430 88 434 92
rect 510 88 514 92
rect 558 88 562 92
rect 598 88 602 92
rect 142 78 146 82
rect 262 78 266 82
rect 294 78 298 82
rect 382 78 386 82
rect 30 68 34 72
rect 78 68 82 72
rect 86 68 90 72
rect 110 68 114 72
rect 142 68 146 72
rect 222 68 226 72
rect 358 68 362 72
rect 542 78 546 82
rect 414 68 418 72
rect 430 68 434 72
rect 526 68 530 72
rect 574 68 578 72
rect 630 68 634 72
rect 158 58 162 62
rect 294 58 298 62
rect 390 58 394 62
rect 406 58 410 62
rect 494 58 498 62
rect 566 58 570 62
rect 102 48 106 52
rect 334 48 338 52
rect 366 48 370 52
rect 6 38 10 42
rect 270 18 274 22
rect 164 3 168 7
rect 169 3 173 7
rect 174 3 178 7
rect 179 3 183 7
rect 184 3 188 7
<< metal2 >>
rect 142 338 146 342
rect 198 338 202 342
rect 214 338 218 342
rect 278 338 282 342
rect 318 338 322 342
rect 414 338 418 342
rect 438 338 442 342
rect 598 341 602 342
rect 598 338 609 341
rect 78 272 81 288
rect 86 272 89 308
rect 106 288 110 291
rect 142 282 145 338
rect 198 312 201 338
rect 158 282 161 308
rect 214 302 217 338
rect 198 292 201 298
rect 278 282 281 338
rect 318 282 321 338
rect 414 282 417 338
rect 378 278 382 281
rect 222 272 225 278
rect 270 272 273 278
rect 278 272 281 278
rect 398 272 401 278
rect 414 272 417 278
rect 438 272 441 338
rect 469 307 475 308
rect 464 303 465 307
rect 469 303 470 307
rect 474 303 475 307
rect 479 303 480 307
rect 469 302 475 303
rect 606 292 609 338
rect 486 272 489 278
rect 346 268 350 271
rect 582 271 585 278
rect 582 268 593 271
rect 18 258 22 261
rect 30 252 33 268
rect 294 262 297 268
rect 518 262 521 268
rect 458 258 462 261
rect 538 258 542 261
rect 54 252 57 258
rect 6 242 9 248
rect 142 162 145 238
rect 186 218 190 221
rect 173 207 179 208
rect 168 203 169 207
rect 173 203 174 207
rect 178 203 179 207
rect 183 203 184 207
rect 173 202 179 203
rect 54 142 57 158
rect 78 152 81 158
rect 134 152 137 158
rect 142 152 145 158
rect 90 148 94 151
rect 186 148 190 151
rect 206 142 209 218
rect 58 138 62 141
rect 162 138 166 141
rect 6 132 9 138
rect 78 132 81 138
rect 94 132 97 138
rect 206 132 209 138
rect 66 128 70 131
rect 106 128 110 131
rect 134 122 137 128
rect 106 118 110 121
rect 30 72 33 118
rect 86 72 89 78
rect 106 68 110 71
rect 134 71 137 118
rect 142 82 145 88
rect 134 68 142 71
rect 78 62 81 68
rect 150 61 153 118
rect 198 92 201 118
rect 214 92 217 258
rect 250 218 254 221
rect 222 162 225 168
rect 266 158 270 161
rect 230 132 233 158
rect 278 142 281 218
rect 302 152 305 218
rect 334 162 337 258
rect 358 252 361 258
rect 414 252 417 258
rect 386 248 390 251
rect 334 142 337 158
rect 358 142 361 218
rect 398 161 401 238
rect 566 192 569 268
rect 582 252 585 258
rect 426 168 430 171
rect 454 162 457 168
rect 398 158 406 161
rect 426 158 430 161
rect 390 152 393 158
rect 406 152 409 158
rect 430 142 433 148
rect 534 142 537 188
rect 574 172 577 218
rect 590 182 593 268
rect 594 158 598 161
rect 394 138 398 141
rect 450 138 454 141
rect 474 138 478 141
rect 530 138 534 141
rect 326 132 329 138
rect 358 132 361 138
rect 542 132 545 158
rect 614 152 617 258
rect 646 242 649 248
rect 622 152 625 158
rect 386 128 390 131
rect 238 122 241 128
rect 226 88 230 91
rect 262 82 265 118
rect 294 82 297 88
rect 222 72 225 78
rect 226 68 230 71
rect 302 71 305 118
rect 294 68 305 71
rect 294 62 297 68
rect 150 58 158 61
rect 150 52 153 58
rect 334 52 337 118
rect 358 72 361 78
rect 366 52 369 118
rect 430 92 433 128
rect 458 118 462 121
rect 469 107 475 108
rect 464 103 465 107
rect 469 103 470 107
rect 474 103 475 107
rect 479 103 480 107
rect 469 102 475 103
rect 502 92 505 128
rect 510 92 513 118
rect 558 92 561 138
rect 566 122 569 138
rect 614 132 617 138
rect 402 88 406 91
rect 602 88 606 91
rect 386 78 390 81
rect 526 72 529 78
rect 542 72 545 78
rect 630 72 633 178
rect 646 142 649 148
rect 410 68 414 71
rect 570 68 574 71
rect 390 62 393 68
rect 430 62 433 68
rect 410 58 414 61
rect 106 48 110 51
rect 6 42 9 48
rect 173 7 179 8
rect 168 3 169 7
rect 173 3 174 7
rect 178 3 179 7
rect 183 3 184 7
rect 173 2 179 3
rect 270 -19 273 18
rect 494 -18 497 58
rect 526 12 529 68
rect 562 58 566 61
rect 574 12 577 68
rect 510 -18 513 8
rect 590 -18 593 8
rect 278 -19 282 -18
rect 270 -22 282 -19
rect 494 -22 498 -18
rect 510 -22 514 -18
rect 590 -22 594 -18
<< m3contact >>
rect 86 308 90 312
rect 78 288 82 292
rect 110 288 114 292
rect 158 308 162 312
rect 198 308 202 312
rect 198 298 202 302
rect 214 298 218 302
rect 222 278 226 282
rect 270 278 274 282
rect 318 278 322 282
rect 382 278 386 282
rect 398 278 402 282
rect 460 303 464 307
rect 465 303 469 307
rect 470 303 474 307
rect 475 303 479 307
rect 480 303 484 307
rect 486 278 490 282
rect 278 268 282 272
rect 294 268 298 272
rect 342 268 346 272
rect 414 268 418 272
rect 14 258 18 262
rect 462 258 466 262
rect 518 258 522 262
rect 534 258 538 262
rect 6 248 10 252
rect 30 248 34 252
rect 54 248 58 252
rect 190 218 194 222
rect 206 218 210 222
rect 164 203 168 207
rect 169 203 173 207
rect 174 203 178 207
rect 179 203 183 207
rect 184 203 188 207
rect 54 158 58 162
rect 78 148 82 152
rect 86 148 90 152
rect 134 148 138 152
rect 142 148 146 152
rect 182 148 186 152
rect 6 138 10 142
rect 62 138 66 142
rect 78 138 82 142
rect 166 138 170 142
rect 206 138 210 142
rect 6 128 10 132
rect 70 128 74 132
rect 94 128 98 132
rect 102 128 106 132
rect 134 128 138 132
rect 110 118 114 122
rect 86 78 90 82
rect 102 68 106 72
rect 142 88 146 92
rect 78 58 82 62
rect 246 218 250 222
rect 278 218 282 222
rect 222 168 226 172
rect 262 158 266 162
rect 358 248 362 252
rect 390 248 394 252
rect 414 248 418 252
rect 302 148 306 152
rect 582 258 586 262
rect 534 188 538 192
rect 566 188 570 192
rect 430 168 434 172
rect 454 168 458 172
rect 406 158 410 162
rect 422 158 426 162
rect 390 148 394 152
rect 430 148 434 152
rect 590 178 594 182
rect 574 168 578 172
rect 598 158 602 162
rect 334 138 338 142
rect 390 138 394 142
rect 454 138 458 142
rect 478 138 482 142
rect 526 138 530 142
rect 646 248 650 252
rect 630 178 634 182
rect 622 158 626 162
rect 614 148 618 152
rect 558 138 562 142
rect 230 128 234 132
rect 326 128 330 132
rect 390 128 394 132
rect 430 128 434 132
rect 542 128 546 132
rect 238 118 242 122
rect 366 118 370 122
rect 198 88 202 92
rect 214 88 218 92
rect 222 88 226 92
rect 294 88 298 92
rect 222 78 226 82
rect 230 68 234 72
rect 358 78 362 82
rect 462 118 466 122
rect 460 103 464 107
rect 465 103 469 107
rect 470 103 474 107
rect 475 103 479 107
rect 480 103 484 107
rect 510 118 514 122
rect 614 128 618 132
rect 566 118 570 122
rect 406 88 410 92
rect 502 88 506 92
rect 606 88 610 92
rect 390 78 394 82
rect 526 78 530 82
rect 646 148 650 152
rect 390 68 394 72
rect 406 68 410 72
rect 542 68 546 72
rect 566 68 570 72
rect 414 58 418 62
rect 430 58 434 62
rect 6 48 10 52
rect 110 48 114 52
rect 150 48 154 52
rect 164 3 168 7
rect 169 3 173 7
rect 174 3 178 7
rect 179 3 183 7
rect 184 3 188 7
rect 558 58 562 62
rect 510 8 514 12
rect 526 8 530 12
rect 574 8 578 12
rect 590 8 594 12
<< metal3 >>
rect 90 308 158 311
rect 162 308 198 311
rect 469 307 475 308
rect 469 302 475 303
rect 202 298 214 301
rect 82 288 110 291
rect 274 278 318 281
rect 386 278 398 281
rect 222 271 225 278
rect 222 268 278 271
rect 298 268 342 271
rect 486 271 489 278
rect 418 268 489 271
rect 18 258 57 261
rect 466 258 518 261
rect 538 258 582 261
rect 54 252 57 258
rect -26 251 -22 252
rect -26 248 6 251
rect 34 248 38 251
rect 362 248 390 251
rect 394 248 414 251
rect 670 251 674 252
rect 650 248 674 251
rect 194 218 206 221
rect 250 218 278 221
rect 173 207 179 208
rect 173 202 179 203
rect 538 188 566 191
rect 594 178 630 181
rect 670 181 674 182
rect 634 178 674 181
rect 422 168 430 171
rect 434 168 454 171
rect 570 168 574 171
rect -26 161 -22 162
rect -26 158 54 161
rect 222 161 225 168
rect 222 158 262 161
rect 410 158 422 161
rect 602 158 622 161
rect 82 148 86 151
rect 90 148 134 151
rect 146 148 182 151
rect 298 148 302 151
rect 394 148 430 151
rect 602 148 614 151
rect 670 151 674 152
rect 650 148 674 151
rect -26 141 -22 142
rect -26 138 6 141
rect 66 138 78 141
rect 170 138 206 141
rect 338 138 390 141
rect 458 138 478 141
rect 482 138 526 141
rect 562 138 617 141
rect 614 132 617 138
rect 10 128 70 131
rect 98 128 102 131
rect 138 128 230 131
rect 330 128 390 131
rect 434 128 542 131
rect 102 118 110 121
rect 114 118 238 121
rect 370 118 462 121
rect 514 118 566 121
rect 469 107 475 108
rect 469 102 475 103
rect 146 88 198 91
rect 218 88 222 91
rect 398 88 406 91
rect 410 88 502 91
rect 602 88 606 91
rect 294 82 297 88
rect 34 78 86 81
rect 90 78 222 81
rect 382 78 390 81
rect 394 78 526 81
rect 78 68 102 71
rect 358 71 361 78
rect 234 68 361 71
rect 394 68 406 71
rect 546 68 566 71
rect 78 62 81 68
rect 418 58 430 61
rect 562 58 566 61
rect -26 51 -22 52
rect -26 48 6 51
rect 114 48 150 51
rect 514 8 526 11
rect 578 8 590 11
rect 173 7 179 8
rect 173 2 179 3
<< m4contact >>
rect 461 303 464 307
rect 464 303 465 307
rect 467 303 469 307
rect 469 303 470 307
rect 470 303 471 307
rect 473 303 474 307
rect 474 303 475 307
rect 475 303 477 307
rect 479 303 480 307
rect 480 303 483 307
rect 38 248 42 252
rect 165 203 168 207
rect 168 203 169 207
rect 171 203 173 207
rect 173 203 174 207
rect 174 203 175 207
rect 177 203 178 207
rect 178 203 179 207
rect 179 203 181 207
rect 183 203 184 207
rect 184 203 187 207
rect 566 168 570 172
rect 294 148 298 152
rect 598 148 602 152
rect 461 103 464 107
rect 464 103 465 107
rect 467 103 469 107
rect 469 103 470 107
rect 470 103 471 107
rect 473 103 474 107
rect 474 103 475 107
rect 475 103 477 107
rect 479 103 480 107
rect 480 103 483 107
rect 598 88 602 92
rect 30 78 34 82
rect 294 78 298 82
rect 566 58 570 62
rect 165 3 168 7
rect 168 3 169 7
rect 171 3 173 7
rect 173 3 174 7
rect 174 3 175 7
rect 177 3 178 7
rect 178 3 179 7
rect 179 3 181 7
rect 183 3 184 7
rect 184 3 187 7
<< metal4 >>
rect 469 307 475 308
rect 469 302 475 303
rect 30 248 38 251
rect 30 82 33 248
rect 173 207 179 208
rect 173 202 179 203
rect 294 82 297 148
rect 469 107 475 108
rect 469 102 475 103
rect 566 62 569 168
rect 598 92 601 148
rect 173 7 179 8
rect 173 2 179 3
<< m5contact >>
rect 460 303 461 307
rect 461 303 464 307
rect 465 303 467 307
rect 467 303 469 307
rect 470 303 471 307
rect 471 303 473 307
rect 473 303 474 307
rect 475 303 477 307
rect 477 303 479 307
rect 480 303 483 307
rect 483 303 484 307
rect 164 203 165 207
rect 165 203 168 207
rect 169 203 171 207
rect 171 203 173 207
rect 174 203 175 207
rect 175 203 177 207
rect 177 203 178 207
rect 179 203 181 207
rect 181 203 183 207
rect 184 203 187 207
rect 187 203 188 207
rect 460 103 461 107
rect 461 103 464 107
rect 465 103 467 107
rect 467 103 469 107
rect 470 103 471 107
rect 471 103 473 107
rect 473 103 474 107
rect 475 103 477 107
rect 477 103 479 107
rect 480 103 483 107
rect 483 103 484 107
rect 164 3 165 7
rect 165 3 168 7
rect 169 3 171 7
rect 171 3 173 7
rect 174 3 175 7
rect 175 3 177 7
rect 177 3 178 7
rect 179 3 181 7
rect 181 3 183 7
rect 184 3 187 7
rect 187 3 188 7
<< metal5 >>
rect 469 307 475 308
rect 464 303 465 307
rect 479 303 480 307
rect 471 302 473 303
rect 173 207 179 208
rect 168 203 169 207
rect 183 203 184 207
rect 175 202 177 203
rect 469 107 475 108
rect 464 103 465 107
rect 479 103 480 107
rect 471 102 473 103
rect 173 7 179 8
rect 168 3 169 7
rect 183 3 184 7
rect 175 2 177 3
<< m6contact >>
rect 466 303 469 307
rect 469 303 470 307
rect 470 303 471 307
rect 473 303 474 307
rect 474 303 475 307
rect 475 303 478 307
rect 466 302 471 303
rect 473 302 478 303
rect 170 203 173 207
rect 173 203 174 207
rect 174 203 175 207
rect 177 203 178 207
rect 178 203 179 207
rect 179 203 182 207
rect 170 202 175 203
rect 177 202 182 203
rect 466 103 469 107
rect 469 103 470 107
rect 470 103 471 107
rect 473 103 474 107
rect 474 103 475 107
rect 475 103 478 107
rect 466 102 471 103
rect 473 102 478 103
rect 170 3 173 7
rect 173 3 174 7
rect 174 3 175 7
rect 177 3 178 7
rect 178 3 179 7
rect 179 3 182 7
rect 170 2 175 3
rect 177 2 182 3
<< metal6 >>
rect 164 207 188 307
rect 164 202 170 207
rect 175 202 177 207
rect 182 202 188 207
rect 164 7 188 202
rect 164 2 170 7
rect 175 2 177 7
rect 182 2 188 7
rect 164 -6 188 2
rect 460 302 466 307
rect 471 302 473 307
rect 478 302 484 307
rect 460 107 484 302
rect 460 102 466 107
rect 471 102 473 107
rect 478 102 484 107
rect 460 -6 484 102
use BUFX2  _31_
timestamp 1592523827
transform -1 0 28 0 -1 105
box -2 -3 26 103
use XOR2X1  _89_
timestamp 1592523827
transform -1 0 84 0 -1 105
box -2 -3 58 103
use XOR2X1  _61_
timestamp 1592523827
transform -1 0 60 0 1 105
box -2 -3 58 103
use INVX1  _58_
timestamp 1592523827
transform 1 0 60 0 1 105
box -2 -3 18 103
use NAND2X1  _76_
timestamp 1592523827
transform 1 0 84 0 -1 105
box -2 -3 26 103
use NAND2X1  _77_
timestamp 1592523827
transform -1 0 132 0 -1 105
box -2 -3 26 103
use INVX1  _57_
timestamp 1592523827
transform 1 0 76 0 1 105
box -2 -3 18 103
use NOR2X1  _59_
timestamp 1592523827
transform -1 0 116 0 1 105
box -2 -3 26 103
use NAND2X1  _60_
timestamp 1592523827
transform 1 0 116 0 1 105
box -2 -3 26 103
use INVX1  _75_
timestamp 1592523827
transform -1 0 148 0 -1 105
box -2 -3 18 103
use AND2X2  _81_
timestamp 1592523827
transform 1 0 148 0 -1 105
box -2 -3 34 103
use NAND2X1  _55_
timestamp 1592523827
transform -1 0 164 0 1 105
box -2 -3 26 103
use FILL  SFILL1800x50
timestamp 1592523827
transform -1 0 188 0 -1 105
box -2 -3 10 103
use FILL  SFILL1640x1050
timestamp 1592523827
transform 1 0 164 0 1 105
box -2 -3 10 103
use FILL  SFILL1720x1050
timestamp 1592523827
transform 1 0 172 0 1 105
box -2 -3 10 103
use FILL  SFILL1800x1050
timestamp 1592523827
transform 1 0 180 0 1 105
box -2 -3 10 103
use NAND2X1  _83_
timestamp 1592523827
transform -1 0 228 0 -1 105
box -2 -3 26 103
use NAND2X1  _84_
timestamp 1592523827
transform -1 0 252 0 -1 105
box -2 -3 26 103
use NOR2X1  _54_
timestamp 1592523827
transform -1 0 212 0 1 105
box -2 -3 26 103
use NAND2X1  _79_
timestamp 1592523827
transform 1 0 212 0 1 105
box -2 -3 26 103
use INVX1  _78_
timestamp 1592523827
transform 1 0 236 0 1 105
box -2 -3 18 103
use FILL  SFILL1880x50
timestamp 1592523827
transform -1 0 196 0 -1 105
box -2 -3 10 103
use FILL  SFILL1960x50
timestamp 1592523827
transform -1 0 204 0 -1 105
box -2 -3 10 103
use INVX1  _82_
timestamp 1592523827
transform -1 0 268 0 -1 105
box -2 -3 18 103
use BUFX2  _29_
timestamp 1592523827
transform -1 0 292 0 -1 105
box -2 -3 26 103
use INVX1  _68_
timestamp 1592523827
transform 1 0 292 0 -1 105
box -2 -3 18 103
use NAND2X1  _70_
timestamp 1592523827
transform 1 0 308 0 -1 105
box -2 -3 26 103
use NAND2X1  _80_
timestamp 1592523827
transform 1 0 252 0 1 105
box -2 -3 26 103
use XOR2X1  _87_
timestamp 1592523827
transform -1 0 332 0 1 105
box -2 -3 58 103
use INVX1  _72_
timestamp 1592523827
transform 1 0 332 0 -1 105
box -2 -3 18 103
use NAND2X1  _74_
timestamp 1592523827
transform 1 0 348 0 -1 105
box -2 -3 26 103
use NAND2X1  _69_
timestamp 1592523827
transform -1 0 356 0 1 105
box -2 -3 26 103
use INVX1  _65_
timestamp 1592523827
transform 1 0 356 0 1 105
box -2 -3 18 103
use INVX1  _37_
timestamp 1592523827
transform -1 0 388 0 -1 105
box -2 -3 18 103
use NOR2X1  _39_
timestamp 1592523827
transform 1 0 388 0 -1 105
box -2 -3 26 103
use NAND2X1  _40_
timestamp 1592523827
transform 1 0 412 0 -1 105
box -2 -3 26 103
use NAND2X1  _67_
timestamp 1592523827
transform 1 0 372 0 1 105
box -2 -3 26 103
use AND2X2  _71_
timestamp 1592523827
transform 1 0 396 0 1 105
box -2 -3 34 103
use NAND2X1  _66_
timestamp 1592523827
transform -1 0 452 0 1 105
box -2 -3 26 103
use INVX1  _38_
timestamp 1592523827
transform -1 0 452 0 -1 105
box -2 -3 18 103
use XOR2X1  _41_
timestamp 1592523827
transform -1 0 532 0 -1 105
box -2 -3 58 103
use NAND2X1  _73_
timestamp 1592523827
transform -1 0 476 0 1 105
box -2 -3 26 103
use FILL  SFILL4520x50
timestamp 1592523827
transform -1 0 460 0 -1 105
box -2 -3 10 103
use FILL  SFILL4600x50
timestamp 1592523827
transform -1 0 468 0 -1 105
box -2 -3 10 103
use FILL  SFILL4680x50
timestamp 1592523827
transform -1 0 476 0 -1 105
box -2 -3 10 103
use FILL  SFILL4760x1050
timestamp 1592523827
transform 1 0 476 0 1 105
box -2 -3 10 103
use FILL  SFILL4840x1050
timestamp 1592523827
transform 1 0 484 0 1 105
box -2 -3 10 103
use INVX1  _33_
timestamp 1592523827
transform -1 0 548 0 -1 105
box -2 -3 18 103
use NOR2X1  _35_
timestamp 1592523827
transform 1 0 548 0 -1 105
box -2 -3 26 103
use INVX1  _62_
timestamp 1592523827
transform 1 0 500 0 1 105
box -2 -3 18 103
use NAND2X1  _64_
timestamp 1592523827
transform 1 0 516 0 1 105
box -2 -3 26 103
use NAND2X1  _63_
timestamp 1592523827
transform -1 0 564 0 1 105
box -2 -3 26 103
use FILL  SFILL4920x1050
timestamp 1592523827
transform 1 0 492 0 1 105
box -2 -3 10 103
use XOR2X1  _36_
timestamp 1592523827
transform 1 0 572 0 -1 105
box -2 -3 58 103
use XOR2X1  _85_
timestamp 1592523827
transform -1 0 620 0 1 105
box -2 -3 58 103
use BUFX2  _27_
timestamp 1592523827
transform 1 0 620 0 1 105
box -2 -3 26 103
use FILL  FILL5800x50
timestamp 1592523827
transform -1 0 636 0 -1 105
box -2 -3 10 103
use FILL  FILL5880x50
timestamp 1592523827
transform -1 0 644 0 -1 105
box -2 -3 10 103
use BUFX2  _30_
timestamp 1592523827
transform -1 0 28 0 -1 305
box -2 -3 26 103
use XOR2X1  _88_
timestamp 1592523827
transform 1 0 28 0 -1 305
box -2 -3 58 103
use XOR2X1  _56_
timestamp 1592523827
transform 1 0 84 0 -1 305
box -2 -3 58 103
use INVX1  _53_
timestamp 1592523827
transform 1 0 140 0 -1 305
box -2 -3 18 103
use INVX1  _52_
timestamp 1592523827
transform 1 0 156 0 -1 305
box -2 -3 18 103
use FILL  SFILL1720x2050
timestamp 1592523827
transform -1 0 180 0 -1 305
box -2 -3 10 103
use FILL  SFILL1800x2050
timestamp 1592523827
transform -1 0 188 0 -1 305
box -2 -3 10 103
use BUFX2  _32_
timestamp 1592523827
transform -1 0 220 0 -1 305
box -2 -3 26 103
use XOR2X1  _51_
timestamp 1592523827
transform 1 0 220 0 -1 305
box -2 -3 58 103
use FILL  SFILL1880x2050
timestamp 1592523827
transform -1 0 196 0 -1 305
box -2 -3 10 103
use INVX1  _47_
timestamp 1592523827
transform 1 0 276 0 -1 305
box -2 -3 18 103
use NOR2X1  _49_
timestamp 1592523827
transform 1 0 292 0 -1 305
box -2 -3 26 103
use INVX1  _48_
timestamp 1592523827
transform 1 0 316 0 -1 305
box -2 -3 18 103
use NAND2X1  _50_
timestamp 1592523827
transform -1 0 356 0 -1 305
box -2 -3 26 103
use NOR2X1  _44_
timestamp 1592523827
transform -1 0 380 0 -1 305
box -2 -3 26 103
use NAND2X1  _45_
timestamp 1592523827
transform -1 0 404 0 -1 305
box -2 -3 26 103
use INVX1  _42_
timestamp 1592523827
transform -1 0 420 0 -1 305
box -2 -3 18 103
use INVX1  _43_
timestamp 1592523827
transform -1 0 436 0 -1 305
box -2 -3 18 103
use XOR2X1  _46_
timestamp 1592523827
transform -1 0 492 0 -1 305
box -2 -3 58 103
use XOR2X1  _86_
timestamp 1592523827
transform -1 0 572 0 -1 305
box -2 -3 58 103
use FILL  SFILL4920x2050
timestamp 1592523827
transform -1 0 500 0 -1 305
box -2 -3 10 103
use FILL  SFILL5000x2050
timestamp 1592523827
transform -1 0 508 0 -1 305
box -2 -3 10 103
use FILL  SFILL5080x2050
timestamp 1592523827
transform -1 0 516 0 -1 305
box -2 -3 10 103
use INVX1  _34_
timestamp 1592523827
transform -1 0 588 0 -1 305
box -2 -3 18 103
use BUFX2  _28_
timestamp 1592523827
transform 1 0 588 0 -1 305
box -2 -3 26 103
use BUFX2  _26_
timestamp 1592523827
transform 1 0 612 0 -1 305
box -2 -3 26 103
use FILL  FILL5880x2050
timestamp 1592523827
transform -1 0 644 0 -1 305
box -2 -3 10 103
<< labels >>
flabel metal6 s 460 -6 484 0 7 FreeSans 24 270 0 0 gnd
port 0 nsew
flabel metal6 s 164 -6 188 0 7 FreeSans 24 270 0 0 vdd
port 1 nsew
flabel metal2 s 214 338 218 342 3 FreeSans 24 90 0 0 s[6]
port 2 nsew
flabel metal3 s -26 48 -22 52 7 FreeSans 24 270 0 0 s[5]
port 3 nsew
flabel metal3 s -26 248 -22 252 7 FreeSans 24 90 0 0 s[4]
port 4 nsew
flabel metal2 s 278 -22 282 -18 7 FreeSans 24 270 0 0 s[3]
port 5 nsew
flabel metal2 s 598 338 602 342 3 FreeSans 24 90 0 0 s[2]
port 6 nsew
flabel metal3 s 670 148 674 152 3 FreeSans 24 0 0 0 s[1]
port 7 nsew
flabel metal3 s 670 248 674 252 3 FreeSans 24 90 0 0 s[0]
port 8 nsew
flabel metal3 s -26 138 -22 142 7 FreeSans 24 0 0 0 x[5]
port 9 nsew
flabel metal2 s 142 338 146 342 3 FreeSans 24 90 0 0 x[4]
port 10 nsew
flabel metal2 s 318 338 322 342 3 FreeSans 24 90 0 0 x[3]
port 11 nsew
flabel metal2 s 438 338 442 342 3 FreeSans 24 90 0 0 x[2]
port 12 nsew
flabel metal2 s 494 -22 498 -18 7 FreeSans 24 270 0 0 x[1]
port 13 nsew
flabel metal3 s 670 178 674 182 3 FreeSans 24 0 0 0 x[0]
port 14 nsew
flabel metal3 s -26 158 -22 162 7 FreeSans 24 0 0 0 y[5]
port 15 nsew
flabel metal2 s 198 338 202 342 3 FreeSans 24 90 0 0 y[4]
port 16 nsew
flabel metal2 s 278 338 282 342 3 FreeSans 24 90 0 0 y[3]
port 17 nsew
flabel metal2 s 414 338 418 342 3 FreeSans 24 90 0 0 y[2]
port 18 nsew
flabel metal2 s 510 -22 514 -18 7 FreeSans 24 270 0 0 y[1]
port 19 nsew
flabel metal2 s 590 -22 594 -18 3 FreeSans 24 270 0 0 y[0]
port 20 nsew
<< end >>
